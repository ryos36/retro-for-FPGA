module retro_main
  (
    input wire clk,
    input wire rst,
    input wire retro_main_ready,
    input wire retro_main_accept,
    output reg retro_main_valid,
    input wire signed [31:0] retro_main_in_memory_q,
    input wire [14:0] retro_main_in_memory_len,
    output wire signed [14:0] retro_main_in_memory_addr,
    output wire signed [31:0] retro_main_in_memory_d,
    output wire retro_main_in_memory_we,
    output wire retro_main_in_memory_req,
    input wire signed [31:0] retro_main_in_io_ports_q,
    input wire [4:0] retro_main_in_io_ports_len,
    output wire signed [4:0] retro_main_in_io_ports_addr,
    output wire signed [31:0] retro_main_in_io_ports_d,
    output wire retro_main_in_io_ports_we,
    output wire retro_main_in_io_ports_req
  );

  //localparams
  localparam retro_main_b1_INIT = 0;
  localparam retro_main_b1_S0 = 1;
  localparam retro_main_b1_S1 = 2;
  localparam retro_main_b1_S2 = 3;
  localparam retro_main_b1_S3 = 4;
  localparam retro_main_b1_S4 = 5;
  localparam retro_main_b1_S5 = 6;
  localparam retro_main_b1_S6 = 7;
  localparam retro_main_b1_S7 = 8;
  localparam retro_main_b1_S8 = 9;
  localparam retro_main_b1_S9 = 10;
  localparam retro_main_b1_S10 = 11;
  localparam retro_main_b1_S11 = 12;
  localparam retro_main_b1_S12 = 13;
  localparam retro_main_b1_S13 = 14;
  localparam retro_main_b1_S14 = 15;
  localparam retro_main_b1_S15 = 16;
  localparam retro_main_b1_S16 = 17;
  localparam retro_main_b1_S17 = 18;
  localparam retro_main_b1_S18 = 19;
  localparam retro_main_b1_S19 = 20;
  localparam retro_main_b1_S20 = 21;
  localparam retro_main_b1_S21 = 22;
  localparam retro_main_b1_S22 = 23;
  localparam retro_main_b1_S23 = 24;
  localparam retro_main_b1_S24 = 25;
  localparam retro_main_b1_S25 = 26;
  localparam retro_main_b1_S26 = 27;
  localparam retro_main_b1_S27 = 28;
  localparam retro_main_b1_S28 = 29;
  localparam retro_main_b1_S29 = 30;
  localparam retro_main_b1_S30 = 31;
  localparam retro_main_b1_S31 = 32;
  localparam retro_main_b1_S32 = 33;
  localparam retro_main_b1_S33 = 34;
  localparam retro_main_b1_S34 = 35;
  localparam retro_main_b1_S35 = 36;
  localparam retro_main_b1_S36 = 37;
  localparam retro_main_b1_S37 = 38;
  localparam retro_main_b1_S38 = 39;
  localparam retro_main_b1_S39 = 40;
  localparam retro_main_b1_S40 = 41;
  localparam retro_main_b1_S41 = 42;
  localparam retro_main_b1_S42 = 43;
  localparam retro_main_b1_S43 = 44;
  localparam retro_main_b1_S44 = 45;
  localparam retro_main_b1_S45 = 46;
  localparam retro_main_b1_S46 = 47;
  localparam retro_main_b1_S47 = 48;
  localparam retro_main_b1_S48 = 49;
  localparam retro_main_b1_S49 = 50;
  localparam retro_main_b1_S50 = 51;
  localparam retro_main_b1_S51 = 52;
  localparam retro_main_b1_S52 = 53;
  localparam retro_main_b1_S53 = 54;
  localparam retro_main_b1_S54 = 55;
  localparam retro_main_b1_S55 = 56;
  localparam retro_main_b1_S56 = 57;
  localparam retro_main_b1_S57 = 58;
  localparam retro_main_b1_S58 = 59;
  localparam retro_main_b1_S59 = 60;
  localparam retro_main_b1_S60 = 61;
  localparam retro_main_b1_S61 = 62;
  localparam retro_main_b1_S62 = 63;
  localparam retro_main_b1_S63 = 64;
  localparam retro_main_b1_S64 = 65;
  localparam retro_main_b1_S65 = 66;
  localparam retro_main_b1_S66 = 67;
  localparam retro_main_b1_S67 = 68;
  localparam retro_main_b1_S68 = 69;
  localparam retro_main_b1_S69 = 70;
  localparam retro_main_b1_S70 = 71;
  localparam retro_main_b1_S71 = 72;
  localparam retro_main_b1_S72 = 73;
  localparam retro_main_b1_S73 = 74;
  localparam retro_main_b1_S74 = 75;
  localparam retro_main_b1_S75 = 76;
  localparam retro_main_b1_S76 = 77;
  localparam retro_main_b1_S77 = 78;
  localparam retro_main_b1_S78 = 79;
  localparam retro_main_b1_S79 = 80;
  localparam retro_main_b1_S80 = 81;
  localparam retro_main_b1_S81 = 82;
  localparam retro_main_b1_S82 = 83;
  localparam retro_main_b1_S83 = 84;
  localparam retro_main_b1_S84 = 85;
  localparam retro_main_b1_S85 = 86;
  localparam retro_main_b1_S86 = 87;
  localparam retro_main_b1_S87 = 88;
  localparam retro_main_b1_S88 = 89;
  localparam retro_main_b1_S89 = 90;
  localparam retro_main_b1_S90 = 91;
  localparam retro_main_b1_S91 = 92;
  localparam retro_main_b1_S92 = 93;
  localparam retro_main_b1_S93 = 94;
  localparam retro_main_b1_S94 = 95;
  localparam retro_main_b1_S95 = 96;
  localparam retro_main_b1_S96 = 97;
  localparam retro_main_b1_S97 = 98;
  localparam retro_main_b1_S98 = 99;
  localparam retro_main_b1_S99 = 100;
  localparam retro_main_b1_S100 = 101;
  localparam retro_main_b1_S101 = 102;
  localparam retro_main_b1_S102 = 103;
  localparam retro_main_b1_S103 = 104;
  localparam retro_main_b1_S104 = 105;
  localparam retro_main_b1_S105 = 106;
  localparam retro_main_b1_S106 = 107;
  localparam retro_main_b1_S107 = 108;
  localparam retro_main_b1_S108 = 109;
  localparam retro_main_b1_S109 = 110;
  localparam retro_main_b1_S110 = 111;
  localparam retro_main_b1_S111 = 112;
  localparam retro_main_b1_S112 = 113;
  localparam retro_main_b1_S113 = 114;
  localparam retro_main_b1_S114 = 115;
  localparam retro_main_b1_S115 = 116;
  localparam retro_main_b1_S116 = 117;
  localparam retro_main_b1_S117 = 118;
  localparam retro_main_b1_S118 = 119;
  localparam retro_main_b1_S119 = 120;
  localparam retro_main_b1_S120 = 121;
  localparam retro_main_b1_S121 = 122;
  localparam retro_main_b1_S122 = 123;
  localparam retro_main_b1_S123 = 124;
  localparam retro_main_b1_S124 = 125;
  localparam retro_main_b1_S125 = 126;
  localparam retro_main_b1_S126 = 127;
  localparam retro_main_b1_S127 = 128;
  localparam retro_main_b1_S128 = 129;
  localparam retro_main_b1_S129 = 130;
  localparam retro_main_b1_S130 = 131;
  localparam retro_main_b1_S131 = 132;
  localparam retro_main_b1_S132 = 133;
  localparam retro_main_b1_S133 = 134;
  localparam retro_main_b1_S134 = 135;
  localparam retro_main_b1_S135 = 136;
  localparam retro_main_b1_S136 = 137;
  localparam retro_main_b1_S137 = 138;
  localparam retro_main_b1_S138 = 139;
  localparam retro_main_b1_S139 = 140;
  localparam retro_main_b1_S140 = 141;
  localparam retro_main_b1_S141 = 142;
  localparam retro_main_b1_S142 = 143;
  localparam retro_main_b1_S143 = 144;
  localparam retro_main_b1_S144 = 145;
  localparam retro_main_b1_S145 = 146;
  localparam retro_main_b1_S146 = 147;
  localparam retro_main_b1_S147 = 148;
  localparam retro_main_b1_S148 = 149;
  localparam retro_main_b1_S149 = 150;
  localparam retro_main_b1_S150 = 151;
  localparam retro_main_b1_S151 = 152;
  localparam retro_main_b1_S152 = 153;
  localparam retro_main_b1_S153 = 154;
  localparam retro_main_b1_S154 = 155;
  localparam retro_main_b1_S155 = 156;
  localparam retro_main_b1_S156 = 157;
  localparam retro_main_b1_S157 = 158;
  localparam retro_main_b1_S158 = 159;
  localparam retro_main_b1_S159 = 160;
  localparam retro_main_b1_S160 = 161;
  localparam retro_main_b1_S161 = 162;
  localparam retro_main_b1_S162 = 163;
  localparam retro_main_b1_S163 = 164;
  localparam retro_main_b1_S164 = 165;
  localparam retro_main_b1_S165 = 166;
  localparam retro_main_b1_S166 = 167;
  localparam retro_main_b1_S167 = 168;
  localparam retro_main_b1_S168 = 169;
  localparam retro_main_b1_S169 = 170;
  localparam retro_main_b1_S170 = 171;
  localparam retro_main_b1_S171 = 172;
  localparam retro_main_b1_S172 = 173;
  localparam retro_main_b1_S173 = 174;
  localparam retro_main_b1_S174 = 175;
  localparam retro_main_b1_S175 = 176;
  localparam retro_main_b1_S176 = 177;
  localparam retro_main_b1_S177 = 178;
  localparam retro_main_b1_S178 = 179;
  localparam retro_main_b1_S179 = 180;
  localparam retro_main_b1_S180 = 181;
  localparam retro_main_b1_S181 = 182;
  localparam retro_main_b1_S182 = 183;
  localparam retro_main_b1_S183 = 184;
  localparam retro_main_b1_S184 = 185;
  localparam retro_main_b1_S185 = 186;
  localparam retro_main_b1_S186 = 187;
  localparam retro_main_b1_S187 = 188;
  localparam retro_main_b1_S188 = 189;
  localparam retro_main_b1_S189 = 190;
  localparam retro_main_b1_S190 = 191;
  localparam retro_main_b1_S191 = 192;
  localparam retro_main_b1_S192 = 193;
  localparam retro_main_b1_S193 = 194;
  localparam retro_main_b1_S194 = 195;
  localparam retro_main_b1_S195 = 196;
  localparam retro_main_b1_S196 = 197;
  localparam retro_main_b1_S197 = 198;
  localparam retro_main_b1_S198 = 199;
  localparam retro_main_b1_S199 = 200;
  localparam retro_main_b1_S200 = 201;
  localparam retro_main_b1_S201 = 202;
  localparam retro_main_b1_S202 = 203;
  localparam retro_main_b1_S203 = 204;
  localparam retro_main_b1_S204 = 205;
  localparam retro_main_b1_S205 = 206;
  localparam retro_main_b1_S206 = 207;
  localparam retro_main_b1_S207 = 208;
  localparam retro_main_b1_S208 = 209;
  localparam retro_main_b1_S209 = 210;
  localparam retro_main_b1_S210 = 211;
  localparam retro_main_b1_S211 = 212;
  localparam retro_main_b1_S212 = 213;
  localparam retro_main_b1_S213 = 214;
  localparam retro_main_b1_S214 = 215;
  localparam retro_main_b1_S215 = 216;
  localparam retro_main_b1_S216 = 217;
  localparam retro_main_b1_S217 = 218;
  localparam retro_main_b1_S218 = 219;
  localparam retro_main_b1_S219 = 220;
  localparam retro_main_b1_S220 = 221;
  localparam retro_main_b1_S221 = 222;
  localparam retro_main_b1_S222 = 223;
  localparam retro_main_b1_S223 = 224;
  localparam retro_main_b1_S224 = 225;
  localparam retro_main_b1_S225 = 226;
  localparam retro_main_b1_S226 = 227;
  localparam retro_main_b1_S227 = 228;
  localparam retro_main_b1_S228 = 229;
  localparam retro_main_b1_S229 = 230;
  localparam retro_main_b1_S230 = 231;
  localparam retro_main_b1_S231 = 232;
  localparam retro_main_b1_S232 = 233;
  localparam retro_main_b1_S233 = 234;
  localparam retro_main_b1_S234 = 235;
  localparam retro_main_b1_S235 = 236;
  localparam retro_main_b1_S236 = 237;
  localparam retro_main_b1_S237 = 238;
  localparam retro_main_b1_S238 = 239;
  localparam retro_main_b1_S239 = 240;
  localparam retro_main_b1_S240 = 241;
  localparam retro_main_b1_S241 = 242;
  localparam retro_main_b1_S242 = 243;
  localparam retro_main_b1_S243 = 244;
  localparam retro_main_b1_S244 = 245;
  localparam retro_main_b1_S245 = 246;
  localparam retro_main_b1_S246 = 247;
  localparam retro_main_b1_S247 = 248;
  localparam retro_main_b1_S248 = 249;
  localparam retro_main_b1_S249 = 250;
  localparam retro_main_b1_S250 = 251;
  localparam retro_main_b1_S251 = 252;
  localparam retro_main_b1_S252 = 253;
  localparam retro_main_b1_S253 = 254;
  localparam retro_main_b1_S254 = 255;
  localparam retro_main_b1_S255 = 256;
  localparam retro_main_b1_S256 = 257;
  localparam retro_main_b1_S257 = 258;
  localparam retro_main_b1_S258 = 259;
  localparam retro_main_b1_S259 = 260;
  localparam retro_main_b1_S260 = 261;
  localparam retro_main_b1_S261 = 262;
  localparam retro_main_b1_S262 = 263;
  localparam retro_main_b1_S263 = 264;
  localparam retro_main_b1_S264 = 265;
  localparam retro_main_b1_S265 = 266;
  localparam retro_main_b1_S266 = 267;
  localparam retro_main_b1_S267 = 268;
  localparam retro_main_b1_S268 = 269;
  localparam retro_main_b1_S269 = 270;
  localparam retro_main_b1_S270 = 271;
  localparam retro_main_b1_S271 = 272;
  localparam retro_main_b1_S272 = 273;
  localparam retro_main_b1_S273 = 274;
  localparam retro_main_b1_S274 = 275;
  localparam retro_main_b1_S275 = 276;
  localparam retro_main_b1_S276 = 277;
  localparam retro_main_b1_S277 = 278;
  localparam retro_main_b1_S278 = 279;
  localparam retro_main_b1_S279 = 280;
  localparam retro_main_b1_S280 = 281;
  localparam retro_main_b1_S281 = 282;
  localparam retro_main_b1_S282 = 283;
  localparam retro_main_b1_S283 = 284;
  localparam retro_main_b1_S284 = 285;
  localparam retro_main_b1_S285 = 286;
  localparam retro_main_b1_S286 = 287;
  localparam retro_main_b1_S287 = 288;
  localparam retro_main_b1_S288 = 289;
  localparam retro_main_b1_S289 = 290;
  localparam retro_main_b1_S290 = 291;
  localparam retro_main_b1_S291 = 292;
  localparam retro_main_b1_S292 = 293;
  localparam retro_main_b1_S293 = 294;
  localparam retro_main_b1_S294 = 295;
  localparam retro_main_b1_S295 = 296;
  localparam retro_main_b1_S296 = 297;
  localparam retro_main_b1_S297 = 298;
  localparam retro_main_b1_S298 = 299;
  localparam retro_main_b1_S299 = 300;
  localparam retro_main_b1_S300 = 301;
  localparam retro_main_b1_S301 = 302;
  localparam retro_main_b1_S302 = 303;
  localparam retro_main_b1_S303 = 304;
  localparam retro_main_b1_S304 = 305;
  localparam retro_main_b1_S305 = 306;
  localparam retro_main_b1_S306 = 307;
  localparam retro_main_b1_S307 = 308;
  localparam retro_main_b1_S308 = 309;
  localparam retro_main_b1_S309 = 310;
  localparam retro_main_b1_S310 = 311;
  localparam retro_main_b1_S311 = 312;
  localparam retro_main_b1_S312 = 313;
  localparam retro_main_b1_S313 = 314;
  localparam retro_main_b1_S314 = 315;
  localparam retro_main_b1_S315 = 316;
  localparam retro_main_b1_S316 = 317;
  localparam retro_main_b1_S317 = 318;
  localparam retro_main_b1_S318 = 319;
  localparam retro_main_b1_S319 = 320;
  localparam retro_main_b1_S320 = 321;
  localparam retro_main_b1_S321 = 322;
  localparam retro_main_b1_S322 = 323;
  localparam retro_main_b1_S323 = 324;
  localparam retro_main_b1_S324 = 325;
  localparam retro_main_b1_S325 = 326;
  localparam retro_main_b1_S326 = 327;
  localparam retro_main_b1_S327 = 328;
  localparam retro_main_b1_S328 = 329;
  localparam retro_main_b1_S329 = 330;
  localparam retro_main_b1_S330 = 331;
  localparam retro_main_b1_S331 = 332;
  localparam retro_main_b1_S332 = 333;
  localparam retro_main_b1_S333 = 334;
  localparam retro_main_b1_S334 = 335;
  localparam retro_main_b1_S335 = 336;
  localparam retro_main_b1_S336 = 337;
  localparam retro_main_b1_S337 = 338;
  localparam retro_main_b1_S338 = 339;
  localparam retro_main_b1_S339 = 340;
  localparam retro_main_b1_S340 = 341;
  localparam retro_main_b1_S341 = 342;
  localparam retro_main_b1_S342 = 343;
  localparam retro_main_b1_S343 = 344;
  localparam retro_main_b1_S344 = 345;
  localparam retro_main_b1_S345 = 346;
  localparam retro_main_b1_S346 = 347;
  localparam retro_main_b1_S347 = 348;
  localparam retro_main_b1_S348 = 349;
  localparam retro_main_b1_S349 = 350;
  localparam retro_main_b1_S350 = 351;
  localparam retro_main_b1_S351 = 352;
  localparam retro_main_b1_S352 = 353;
  localparam retro_main_b1_S353 = 354;
  localparam retro_main_b1_S354 = 355;
  localparam retro_main_b1_S355 = 356;
  localparam retro_main_b1_S356 = 357;
  localparam retro_main_b1_S357 = 358;
  localparam retro_main_b1_S358 = 359;
  localparam retro_main_b1_S359 = 360;
  localparam retro_main_b1_S360 = 361;
  localparam retro_main_b1_S361 = 362;
  localparam retro_main_b1_S362 = 363;
  localparam retro_main_b1_S363 = 364;
  localparam retro_main_b1_S364 = 365;
  localparam retro_main_b1_S365 = 366;
  localparam retro_main_b1_S366 = 367;
  localparam retro_main_b1_S367 = 368;
  localparam retro_main_b1_S368 = 369;
  localparam retro_main_b1_S369 = 370;
  localparam retro_main_b1_S370 = 371;
  localparam retro_main_b1_S371 = 372;
  localparam retro_main_b1_S372 = 373;
  localparam retro_main_b1_S373 = 374;
  localparam retro_main_b1_S374 = 375;
  localparam retro_main_b1_S375 = 376;
  localparam retro_main_b1_S376 = 377;
  localparam retro_main_b1_S377 = 378;
  localparam retro_main_b1_S378 = 379;
  localparam retro_main_b1_S379 = 380;
  localparam retro_main_b1_S380 = 381;
  localparam retro_main_b1_S381 = 382;
  localparam retro_main_b1_S382 = 383;
  localparam retro_main_b1_S383 = 384;
  localparam retro_main_b1_S384 = 385;
  localparam retro_main_b1_S385 = 386;
  localparam retro_main_b1_S386 = 387;
  localparam retro_main_b1_S387 = 388;
  localparam retro_main_b1_S388 = 389;
  localparam retro_main_b1_S389 = 390;
  localparam retro_main_b1_S390 = 391;
  localparam retro_main_b1_S391 = 392;
  localparam retro_main_b1_S392 = 393;
  localparam retro_main_b1_S393 = 394;
  localparam retro_main_b1_S394 = 395;
  localparam retro_main_b1_S395 = 396;
  localparam retro_main_b1_S396 = 397;
  localparam retro_main_b1_S397 = 398;
  localparam retro_main_b1_S398 = 399;
  localparam retro_main_b1_S399 = 400;
  localparam retro_main_b1_S400 = 401;
  localparam retro_main_b1_S401 = 402;
  localparam retro_main_b1_S402 = 403;
  localparam retro_main_b1_S403 = 404;
  localparam retro_main_b1_S404 = 405;
  localparam retro_main_b1_S405 = 406;
  localparam retro_main_b1_S406 = 407;
  localparam retro_main_b1_S407 = 408;
  localparam retro_main_b1_S408 = 409;
  localparam retro_main_b1_S409 = 410;
  localparam retro_main_b1_S410 = 411;
  localparam retro_main_b1_S411 = 412;
  localparam retro_main_b1_S412 = 413;
  localparam retro_main_b1_S413 = 414;
  localparam retro_main_b1_S414 = 415;
  localparam retro_main_b1_S415 = 416;
  localparam retro_main_b1_S416 = 417;
  localparam retro_main_b1_S417 = 418;
  localparam retro_main_b1_S418 = 419;
  localparam retro_main_b1_S419 = 420;
  localparam retro_main_b1_S420 = 421;
  localparam retro_main_b1_S421 = 422;
  localparam retro_main_b1_S422 = 423;
  localparam retro_main_b1_S423 = 424;
  localparam retro_main_b1_S424 = 425;
  localparam retro_main_b1_S425 = 426;
  localparam retro_main_b1_S426 = 427;
  localparam retro_main_b1_S427 = 428;
  localparam retro_main_b1_S428 = 429;
  localparam retro_main_b1_S429 = 430;
  localparam retro_main_b1_S430 = 431;
  localparam retro_main_b1_S431 = 432;
  localparam retro_main_b1_S432 = 433;
  localparam retro_main_b1_S433 = 434;
  localparam retro_main_b1_S434 = 435;
  localparam retro_main_b1_S435 = 436;
  localparam retro_main_b1_S436 = 437;
  localparam retro_main_b1_S437 = 438;
  localparam retro_main_b1_S438 = 439;
  localparam retro_main_b1_S439 = 440;
  localparam retro_main_b1_S440 = 441;
  localparam retro_main_b1_S441 = 442;
  localparam retro_main_b1_S442 = 443;
  localparam retro_main_b1_S443 = 444;
  localparam retro_main_b1_S444 = 445;
  localparam retro_main_b1_S445 = 446;
  localparam retro_main_b1_S446 = 447;
  localparam retro_main_b1_S447 = 448;
  localparam retro_main_b1_S448 = 449;
  localparam retro_main_b1_S449 = 450;
  localparam retro_main_b1_S450 = 451;
  localparam retro_main_b1_S451 = 452;
  localparam retro_main_b1_S452 = 453;
  localparam retro_main_b1_S453 = 454;
  localparam retro_main_b1_S454 = 455;
  localparam retro_main_b1_S455 = 456;
  localparam retro_main_b1_S456 = 457;
  localparam retro_main_b1_S457 = 458;
  localparam retro_main_b1_S458 = 459;
  localparam retro_main_b1_S459 = 460;
  localparam retro_main_b1_S460 = 461;
  localparam retro_main_b1_S461 = 462;
  localparam retro_main_b1_S462 = 463;
  localparam retro_main_b1_S463 = 464;
  localparam retro_main_b1_S464 = 465;
  localparam retro_main_b1_S465 = 466;
  localparam retro_main_b1_S466 = 467;
  localparam retro_main_b1_S467 = 468;
  localparam retro_main_b1_S468 = 469;
  localparam retro_main_b1_S469 = 470;
  localparam retro_main_b1_S470 = 471;
  localparam retro_main_b1_S471 = 472;
  localparam retro_main_b1_S472 = 473;
  localparam retro_main_b1_S473 = 474;
  localparam retro_main_b1_S474 = 475;
  localparam retro_main_b1_S475 = 476;
  localparam retro_main_b1_S476 = 477;
  localparam retro_main_b1_S477 = 478;
  localparam retro_main_b1_S478 = 479;
  localparam retro_main_b1_S479 = 480;
  localparam retro_main_b1_S480 = 481;
  localparam retro_main_b1_S481 = 482;
  localparam retro_main_b1_S482 = 483;
  localparam retro_main_b1_S483 = 484;
  localparam retro_main_b1_S484 = 485;
  localparam retro_main_b1_S485 = 486;
  localparam retro_main_b1_S486 = 487;
  localparam retro_main_b1_S487 = 488;
  localparam retro_main_b1_S488 = 489;
  localparam retro_main_b1_S489 = 490;
  localparam retro_main_b1_S490 = 491;
  localparam retro_main_b1_S491 = 492;
  localparam retro_main_b1_S492 = 493;
  localparam retro_main_b1_S493 = 494;
  localparam retro_main_b1_S494 = 495;
  localparam retro_main_b1_S495 = 496;
  localparam retro_main_b1_S496 = 497;
  localparam retro_main_b1_S497 = 498;
  localparam retro_main_b1_S498 = 499;
  localparam retro_main_b1_S499 = 500;
  localparam retro_main_b1_S500 = 501;
  localparam retro_main_b1_S501 = 502;
  localparam retro_main_b1_S502 = 503;
  localparam retro_main_b1_S503 = 504;
  localparam retro_main_b1_S504 = 505;
  localparam retro_main_b1_S505 = 506;
  localparam retro_main_b1_S506 = 507;
  localparam retro_main_b1_S507 = 508;
  localparam retro_main_b1_S508 = 509;
  localparam retro_main_b1_S509 = 510;
  localparam retro_main_b1_S510 = 511;
  localparam retro_main_b1_S511 = 512;
  localparam retro_main_b1_S512 = 513;
  localparam retro_main_b1_S513 = 514;
  localparam retro_main_b1_S514 = 515;
  localparam retro_main_b1_S515 = 516;
  localparam retro_main_b1_S516 = 517;
  localparam retro_main_b1_S517 = 518;
  localparam retro_main_b1_S518 = 519;
  localparam retro_main_b1_S519 = 520;
  localparam retro_main_b1_S520 = 521;
  localparam retro_main_b1_S521 = 522;
  localparam retro_main_b1_S522 = 523;
  localparam retro_main_b1_S523 = 524;
  localparam retro_main_b1_S524 = 525;
  localparam retro_main_b1_S525 = 526;
  localparam retro_main_b1_S526 = 527;
  localparam retro_main_b1_S527 = 528;
  localparam retro_main_b1_S528 = 529;
  localparam retro_main_b1_S529 = 530;
  localparam retro_main_b1_S530 = 531;
  localparam retro_main_b1_S531 = 532;
  localparam retro_main_b1_S532 = 533;
  localparam retro_main_b1_S533 = 534;
  localparam retro_main_b1_S534 = 535;
  localparam retro_main_b1_S535 = 536;
  localparam retro_main_b1_S536 = 537;
  localparam retro_main_b1_S537 = 538;
  localparam retro_main_b1_S538 = 539;
  localparam retro_main_b1_S539 = 540;
  localparam retro_main_b1_S540 = 541;
  localparam retro_main_b1_S541 = 542;
  localparam retro_main_b1_S542 = 543;
  localparam retro_main_b1_S543 = 544;
  localparam retro_main_b1_S544 = 545;
  localparam retro_main_b1_S545 = 546;
  localparam retro_main_b1_S546 = 547;
  localparam retro_main_b1_S547 = 548;
  localparam retro_main_b1_S548 = 549;
  localparam retro_main_b1_S549 = 550;
  localparam retro_main_b1_S550 = 551;
  localparam retro_main_b1_S551 = 552;
  localparam retro_main_b1_S552 = 553;
  localparam retro_main_b1_S553 = 554;
  localparam retro_main_b1_S554 = 555;
  localparam retro_main_b1_S555 = 556;
  localparam retro_main_b1_S556 = 557;
  localparam retro_main_b1_S557 = 558;
  localparam retro_main_b1_S558 = 559;
  localparam retro_main_b1_S559 = 560;
  localparam retro_main_b1_S560 = 561;
  localparam retro_main_b1_S561 = 562;
  localparam retro_main_b1_S562 = 563;
  localparam retro_main_b1_S563 = 564;
  localparam retro_main_b1_S564 = 565;
  localparam retro_main_b1_S565 = 566;
  localparam retro_main_b1_S566 = 567;
  localparam retro_main_b1_S567 = 568;
  localparam retro_main_b1_S568 = 569;
  localparam retro_main_b1_S569 = 570;
  localparam retro_main_b1_S570 = 571;
  localparam retro_main_b1_S571 = 572;
  localparam retro_main_b1_S572 = 573;
  localparam retro_main_b1_S573 = 574;
  localparam retro_main_b1_S574 = 575;
  localparam retro_main_b1_S575 = 576;
  localparam retro_main_b1_S576 = 577;
  localparam retro_main_b1_S577 = 578;
  localparam retro_main_b1_S578 = 579;
  localparam retro_main_b1_S579 = 580;
  localparam retro_main_b1_S580 = 581;
  localparam retro_main_b1_S581 = 582;
  localparam retro_main_b1_S582 = 583;
  localparam retro_main_b1_S583 = 584;
  localparam retro_main_b1_S584 = 585;
  localparam retro_main_b1_S585 = 586;
  localparam retro_main_b1_S586 = 587;
  localparam retro_main_b1_S587 = 588;
  localparam retro_main_b1_S588 = 589;
  localparam retro_main_b1_S589 = 590;
  localparam retro_main_b1_S590 = 591;
  localparam retro_main_b1_S591 = 592;
  localparam retro_main_b1_S592 = 593;
  localparam retro_main_b1_S593 = 594;
  localparam retro_main_b1_S594 = 595;
  localparam retro_main_b1_S595 = 596;
  localparam retro_main_b1_S596 = 597;
  localparam retro_main_b1_S597 = 598;
  localparam retro_main_b1_S598 = 599;
  localparam retro_main_b1_S599 = 600;
  localparam retro_main_b1_S600 = 601;
  localparam retro_main_b1_S601 = 602;
  localparam retro_main_b1_S602 = 603;
  localparam retro_main_b1_S603 = 604;
  localparam retro_main_b1_S604 = 605;
  localparam retro_main_b1_S605 = 606;
  localparam retro_main_b1_S606 = 607;
  localparam retro_main_b1_S607 = 608;
  localparam retro_main_b1_S608 = 609;
  localparam retro_main_b1_S609 = 610;
  localparam retro_main_b1_S610 = 611;
  localparam retro_main_b1_S611 = 612;
  localparam retro_main_b1_S612 = 613;
  localparam retro_main_b1_S613 = 614;
  localparam retro_main_b1_S614 = 615;
  localparam retro_main_b1_S615 = 616;
  localparam retro_main_b1_S616 = 617;
  localparam retro_main_b1_S617 = 618;
  localparam retro_main_b1_S618 = 619;
  localparam retro_main_b1_S619 = 620;
  localparam retro_main_b1_S620 = 621;
  localparam retro_main_b1_S621 = 622;
  localparam retro_main_b1_S622 = 623;
  localparam retro_main_b1_S623 = 624;
  localparam retro_main_b1_S624 = 625;
  localparam retro_main_b1_S625 = 626;
  localparam retro_main_b1_S626 = 627;
  localparam retro_main_b1_S627 = 628;
  localparam retro_main_b1_S628 = 629;
  localparam retro_main_b1_S629 = 630;
  localparam retro_main_b1_S630 = 631;
  localparam retro_main_b1_S631 = 632;
  localparam retro_main_b1_S632 = 633;
  localparam retro_main_b1_S633 = 634;
  localparam retro_main_b1_S634 = 635;
  localparam retro_main_b1_S635 = 636;
  localparam retro_main_b1_S636 = 637;
  localparam retro_main_b1_S637 = 638;
  localparam retro_main_b1_S638 = 639;
  localparam retro_main_b1_S639 = 640;
  localparam retro_main_b1_S640 = 641;
  localparam retro_main_b1_S641 = 642;
  localparam retro_main_b1_S642 = 643;
  localparam retro_main_b1_S643 = 644;
  localparam retro_main_b1_S644 = 645;
  localparam retro_main_b1_S645 = 646;
  localparam retro_main_b1_S646 = 647;
  localparam retro_main_b1_S647 = 648;
  localparam retro_main_b1_S648 = 649;
  localparam retro_main_b1_S649 = 650;
  localparam retro_main_b1_S650 = 651;
  localparam retro_main_b1_S651 = 652;
  localparam retro_main_b1_S652 = 653;
  localparam retro_main_b1_S653 = 654;
  localparam retro_main_b1_S654 = 655;
  localparam retro_main_b1_S655 = 656;
  localparam retro_main_b1_S656 = 657;
  localparam retro_main_b1_S657 = 658;
  localparam retro_main_b1_S658 = 659;
  localparam retro_main_b1_S659 = 660;
  localparam retro_main_b1_S660 = 661;
  localparam retro_main_b1_S661 = 662;
  localparam retro_main_b1_S662 = 663;
  localparam retro_main_b1_S663 = 664;
  localparam retro_main_b1_S664 = 665;
  localparam retro_main_b1_S665 = 666;
  localparam retro_main_b1_S666 = 667;
  localparam retro_main_b1_S667 = 668;
  localparam retro_main_b1_S668 = 669;
  localparam retro_main_b1_S669 = 670;
  localparam retro_main_b1_S670 = 671;
  localparam retro_main_b1_S671 = 672;
  localparam retro_main_b1_S672 = 673;
  localparam retro_main_b1_S673 = 674;
  localparam retro_main_b1_S674 = 675;
  localparam retro_main_b1_S675 = 676;
  localparam retro_main_b1_S676 = 677;
  localparam retro_main_b1_S677 = 678;
  localparam retro_main_b1_S678 = 679;
  localparam retro_main_b1_S679 = 680;
  localparam retro_main_b1_S680 = 681;
  localparam retro_main_b1_S681 = 682;
  localparam retro_main_b1_S682 = 683;
  localparam retro_main_b1_S683 = 684;
  localparam retro_main_b1_S684 = 685;
  localparam retro_main_b1_S685 = 686;
  localparam retro_main_b1_S686 = 687;
  localparam retro_main_b1_S687 = 688;
  localparam retro_main_b1_S688 = 689;
  localparam retro_main_b1_S689 = 690;
  localparam retro_main_b1_S690 = 691;
  localparam retro_main_b1_S691 = 692;
  localparam retro_main_b1_S692 = 693;
  localparam retro_main_b1_S693 = 694;
  localparam retro_main_b1_S694 = 695;
  localparam retro_main_b1_S695 = 696;
  localparam retro_main_b1_S696 = 697;
  localparam retro_main_b1_S697 = 698;
  localparam retro_main_b1_S698 = 699;
  localparam retro_main_b1_S699 = 700;
  localparam retro_main_b1_S700 = 701;
  localparam retro_main_b1_S701 = 702;
  localparam retro_main_b1_S702 = 703;
  localparam retro_main_b1_S703 = 704;
  localparam retro_main_b1_S704 = 705;
  localparam retro_main_b1_S705 = 706;
  localparam retro_main_b1_S706 = 707;
  localparam retro_main_b1_S707 = 708;
  localparam retro_main_b1_S708 = 709;
  localparam retro_main_b1_S709 = 710;
  localparam retro_main_b1_S710 = 711;
  localparam retro_main_b1_S711 = 712;
  localparam retro_main_b1_S712 = 713;
  localparam retro_main_b1_S713 = 714;
  localparam retro_main_b1_S714 = 715;
  localparam retro_main_b1_S715 = 716;
  localparam retro_main_b1_S716 = 717;
  localparam retro_main_b1_S717 = 718;
  localparam retro_main_b1_S718 = 719;
  localparam retro_main_b1_S719 = 720;
  localparam retro_main_b1_S720 = 721;
  localparam retro_main_b1_S721 = 722;
  localparam retro_main_b1_S722 = 723;
  localparam retro_main_b1_S723 = 724;
  localparam retro_main_b1_S724 = 725;
  localparam retro_main_b1_S725 = 726;
  localparam retro_main_b1_S726 = 727;
  localparam retro_main_b1_S727 = 728;
  localparam retro_main_b1_S728 = 729;
  localparam retro_main_b1_S729 = 730;
  localparam retro_main_b1_S730 = 731;
  localparam retro_main_b1_S731 = 732;
  localparam retro_main_b1_S732 = 733;
  localparam retro_main_b1_S733 = 734;
  localparam retro_main_b1_S734 = 735;
  localparam retro_main_b1_S735 = 736;
  localparam retro_main_b1_S736 = 737;
  localparam retro_main_b1_S737 = 738;
  localparam retro_main_b1_S738 = 739;
  localparam retro_main_b1_S739 = 740;
  localparam retro_main_b1_S740 = 741;
  localparam retro_main_b1_S741 = 742;
  localparam retro_main_b1_S742 = 743;
  localparam retro_main_b1_S743 = 744;
  localparam retro_main_b1_S744 = 745;
  localparam retro_main_b1_S745 = 746;
  localparam retro_main_b1_S746 = 747;
  localparam retro_main_b1_S747 = 748;
  localparam retro_main_b1_S748 = 749;
  localparam retro_main_b1_S749 = 750;
  localparam retro_main_b1_S750 = 751;
  localparam retro_main_b1_S751 = 752;
  localparam retro_main_b1_S752 = 753;
  localparam retro_main_b1_S753 = 754;
  localparam retro_main_b1_S754 = 755;
  localparam retro_main_b1_S755 = 756;
  localparam retro_main_b1_S756 = 757;
  localparam retro_main_b1_S757 = 758;
  localparam retro_main_b1_S758 = 759;
  localparam retro_main_b1_S759 = 760;
  localparam retro_main_b1_S760 = 761;
  localparam retro_main_b1_S761 = 762;
  localparam retro_main_b1_S762 = 763;
  localparam retro_main_b1_S763 = 764;
  localparam retro_main_b1_S764 = 765;
  localparam retro_main_b1_S765 = 766;
  localparam retro_main_b1_S766 = 767;
  localparam retro_main_b1_S767 = 768;
  localparam retro_main_b1_S768 = 769;
  localparam retro_main_b1_S769 = 770;
  localparam retro_main_b1_S770 = 771;
  localparam retro_main_b1_S771 = 772;
  localparam retro_main_b1_S772 = 773;
  localparam retro_main_b1_S773 = 774;
  localparam retro_main_b1_S774 = 775;
  localparam retro_main_b1_S775 = 776;
  localparam retro_main_b1_S776 = 777;
  localparam retro_main_b1_S777 = 778;
  localparam retro_main_b1_S778 = 779;
  localparam retro_main_b1_S779 = 780;
  localparam retro_main_b1_S780 = 781;
  localparam retro_main_b1_S781 = 782;
  localparam retro_main_b1_S782 = 783;
  localparam retro_main_b1_S783 = 784;
  localparam retro_main_b1_S784 = 785;
  localparam retro_main_b1_S785 = 786;
  localparam retro_main_b1_S786 = 787;
  localparam retro_main_b1_S787 = 788;
  localparam retro_main_b1_S788 = 789;
  localparam retro_main_b1_S789 = 790;
  localparam retro_main_b1_S790 = 791;
  localparam retro_main_b1_S791 = 792;
  localparam retro_main_b1_S792 = 793;
  localparam retro_main_b1_S793 = 794;
  localparam retro_main_b1_S794 = 795;
  localparam retro_main_b1_S795 = 796;
  localparam retro_main_b1_S796 = 797;
  localparam retro_main_b1_S797 = 798;
  localparam retro_main_b1_S798 = 799;
  localparam retro_main_b1_S799 = 800;
  localparam retro_main_b1_S800 = 801;
  localparam retro_main_b1_S801 = 802;
  localparam retro_main_b1_S802 = 803;
  localparam retro_main_b1_S803 = 804;
  localparam retro_main_b1_S804 = 805;
  localparam retro_main_b1_S805 = 806;
  localparam retro_main_b1_S806 = 807;
  localparam retro_main_b1_S807 = 808;
  localparam retro_main_b1_S808 = 809;
  localparam retro_main_b1_S809 = 810;
  localparam retro_main_b1_S810 = 811;
  localparam retro_main_b1_S811 = 812;
  localparam retro_main_b1_S812 = 813;
  localparam retro_main_b1_S813 = 814;
  localparam retro_main_b1_S814 = 815;
  localparam retro_main_b1_S815 = 816;
  localparam retro_main_b1_S816 = 817;
  localparam retro_main_b1_S817 = 818;
  localparam retro_main_b1_S818 = 819;
  localparam retro_main_b1_S819 = 820;
  localparam retro_main_b1_S820 = 821;
  localparam retro_main_b1_S821 = 822;
  localparam retro_main_b1_S822 = 823;
  localparam retro_main_b1_S823 = 824;
  localparam retro_main_b1_S824 = 825;
  localparam retro_main_b1_S825 = 826;
  localparam retro_main_b1_S826 = 827;
  localparam retro_main_b1_S827 = 828;
  localparam retro_main_b1_S828 = 829;
  localparam retro_main_b1_S829 = 830;
  localparam retro_main_b1_S830 = 831;
  localparam retro_main_b1_S831 = 832;
  localparam retro_main_b1_S832 = 833;
  localparam retro_main_b1_S833 = 834;
  localparam retro_main_b1_S834 = 835;
  localparam retro_main_b1_S835 = 836;
  localparam retro_main_b1_S836 = 837;
  localparam retro_main_b1_S837 = 838;
  localparam retro_main_b1_S838 = 839;
  localparam retro_main_b1_S839 = 840;
  localparam retro_main_b1_S840 = 841;
  localparam retro_main_b1_S841 = 842;
  localparam retro_main_b1_S842 = 843;
  localparam retro_main_b1_S843 = 844;
  localparam retro_main_b1_S844 = 845;
  localparam retro_main_b1_S845 = 846;
  localparam retro_main_b1_S846 = 847;
  localparam retro_main_b1_S847 = 848;
  localparam retro_main_b1_S848 = 849;
  localparam retro_main_b1_S849 = 850;
  localparam retro_main_b1_S850 = 851;
  localparam retro_main_b1_S851 = 852;
  localparam retro_main_b1_S852 = 853;
  localparam retro_main_b1_S853 = 854;
  localparam retro_main_b1_S854 = 855;
  localparam retro_main_b1_S855 = 856;
  localparam retro_main_b1_S856 = 857;
  localparam retro_main_b1_S857 = 858;
  localparam retro_main_b1_S858 = 859;
  localparam retro_main_b1_S859 = 860;
  localparam retro_main_b1_S860 = 861;
  localparam retro_main_b1_S861 = 862;
  localparam retro_main_b1_S862 = 863;
  localparam retro_main_b1_S863 = 864;
  localparam retro_main_b1_S864 = 865;
  localparam retro_main_b1_S865 = 866;
  localparam retro_main_b1_S866 = 867;
  localparam retro_main_b1_S867 = 868;
  localparam retro_main_b1_S868 = 869;
  localparam retro_main_b1_S869 = 870;
  localparam retro_main_b1_S870 = 871;
  localparam retro_main_b1_S871 = 872;
  localparam retro_main_b1_S872 = 873;
  localparam retro_main_b1_S873 = 874;
  localparam retro_main_b1_S874 = 875;
  localparam retro_main_b1_S875 = 876;
  localparam retro_main_b1_S876 = 877;
  localparam retro_main_b1_S877 = 878;
  localparam retro_main_b1_S878 = 879;
  localparam retro_main_b1_S879 = 880;
  localparam retro_main_b1_S880 = 881;
  localparam retro_main_b1_S881 = 882;
  localparam retro_main_b1_S882 = 883;
  localparam retro_main_b1_S883 = 884;
  localparam retro_main_b1_S884 = 885;
  localparam retro_main_b1_S885 = 886;
  localparam retro_main_b1_S886 = 887;
  localparam retro_main_b1_S887 = 888;
  localparam retro_main_b1_S888 = 889;
  localparam retro_main_b1_S889 = 890;
  localparam retro_main_b1_S890 = 891;
  localparam retro_main_b1_S891 = 892;
  localparam retro_main_b1_S892 = 893;
  localparam retro_main_b1_S893 = 894;
  localparam retro_main_b1_S894 = 895;
  localparam retro_main_b1_S895 = 896;
  localparam retro_main_b1_S896 = 897;
  localparam retro_main_b1_S897 = 898;
  localparam retro_main_b1_S898 = 899;
  localparam retro_main_b1_S899 = 900;
  localparam retro_main_b1_S900 = 901;
  localparam retro_main_b1_S901 = 902;
  localparam retro_main_b1_S902 = 903;
  localparam retro_main_b1_S903 = 904;
  localparam retro_main_b1_S904 = 905;
  localparam retro_main_b1_S905 = 906;
  localparam retro_main_b1_S906 = 907;
  localparam retro_main_b1_S907 = 908;
  localparam retro_main_b1_S908 = 909;
  localparam retro_main_b1_S909 = 910;
  localparam retro_main_b1_S910 = 911;
  localparam retro_main_b1_S911 = 912;
  localparam retro_main_b1_S912 = 913;
  localparam retro_main_b1_S913 = 914;
  localparam retro_main_b1_S914 = 915;
  localparam retro_main_b1_S915 = 916;
  localparam retro_main_b1_S916 = 917;
  localparam retro_main_b1_S917 = 918;
  localparam retro_main_b1_S918 = 919;
  localparam retro_main_b1_S919 = 920;
  localparam retro_main_b1_S920 = 921;
  localparam retro_main_b1_S921 = 922;
  localparam retro_main_b1_S922 = 923;
  localparam retro_main_b1_S923 = 924;
  localparam retro_main_b1_S924 = 925;
  localparam retro_main_b1_S925 = 926;
  localparam retro_main_b1_S926 = 927;
  localparam retro_main_b1_S927 = 928;
  localparam retro_main_b1_S928 = 929;
  localparam retro_main_b1_S929 = 930;
  localparam retro_main_b1_S930 = 931;
  localparam retro_main_b1_S931 = 932;
  localparam retro_main_b1_S932 = 933;
  localparam retro_main_b1_S933 = 934;
  localparam retro_main_b1_S934 = 935;
  localparam retro_main_b1_S935 = 936;
  localparam retro_main_b1_S936 = 937;
  localparam retro_main_b1_S937 = 938;
  localparam retro_main_b1_S938 = 939;
  localparam retro_main_b1_S939 = 940;
  localparam retro_main_b1_S940 = 941;
  localparam retro_main_b1_S941 = 942;
  localparam retro_main_b1_S942 = 943;
  localparam retro_main_b1_S943 = 944;
  localparam retro_main_b1_S944 = 945;
  localparam retro_main_b1_S945 = 946;
  localparam retro_main_b1_S946 = 947;
  localparam retro_main_b1_S947 = 948;
  localparam retro_main_b1_S948 = 949;
  localparam retro_main_b1_S949 = 950;
  localparam retro_main_b1_S950 = 951;
  localparam retro_main_b1_S951 = 952;
  localparam retro_main_b1_S952 = 953;
  localparam retro_main_b1_S953 = 954;
  localparam retro_main_b1_S954 = 955;
  localparam retro_main_b1_S955 = 956;
  localparam retro_main_b1_S956 = 957;
  localparam retro_main_b1_S957 = 958;
  localparam retro_main_b1_S958 = 959;
  localparam retro_main_b1_S959 = 960;
  localparam retro_main_b1_S960 = 961;
  localparam retro_main_b1_S961 = 962;
  localparam retro_main_b1_S962 = 963;
  localparam retro_main_b1_S963 = 964;
  localparam retro_main_b1_S964 = 965;
  localparam retro_main_b1_S965 = 966;
  localparam retro_main_b1_S966 = 967;
  localparam retro_main_b1_S967 = 968;
  localparam retro_main_b1_S968 = 969;
  localparam retro_main_b1_S969 = 970;
  localparam retro_main_b1_S970 = 971;
  localparam retro_main_b1_S971 = 972;
  localparam retro_main_b1_S972 = 973;
  localparam retro_main_b1_S973 = 974;
  localparam retro_main_b1_S974 = 975;
  localparam retro_main_b1_S975 = 976;
  localparam retro_main_b1_S976 = 977;
  localparam retro_main_b1_S977 = 978;
  localparam retro_main_b1_S978 = 979;
  localparam retro_main_b1_S979 = 980;
  localparam retro_main_b1_S980 = 981;
  localparam retro_main_b1_S981 = 982;
  localparam retro_main_b1_S982 = 983;
  localparam retro_main_b1_S983 = 984;
  localparam retro_main_b1_S984 = 985;
  localparam retro_main_b1_S985 = 986;
  localparam retro_main_b1_S986 = 987;
  localparam retro_main_b1_S987 = 988;
  localparam retro_main_b1_S988 = 989;
  localparam retro_main_b1_S989 = 990;
  localparam retro_main_b1_S990 = 991;
  localparam retro_main_b1_S991 = 992;
  localparam retro_main_b1_S992 = 993;
  localparam retro_main_b1_S993 = 994;
  localparam retro_main_b1_S994 = 995;
  localparam retro_main_b1_S995 = 996;
  localparam retro_main_b1_S996 = 997;
  localparam retro_main_b1_S997 = 998;
  localparam retro_main_b1_S998 = 999;
  localparam retro_main_b1_S999 = 1000;
  localparam retro_main_b1_S1000 = 1001;
  localparam retro_main_b1_S1001 = 1002;
  localparam retro_main_b1_S1002 = 1003;
  localparam retro_main_b1_S1003 = 1004;
  localparam retro_main_b1_S1004 = 1005;
  localparam retro_main_b1_S1005 = 1006;
  localparam retro_main_b1_S1006 = 1007;
  localparam retro_main_b1_S1007 = 1008;
  localparam retro_main_b1_S1008 = 1009;
  localparam retro_main_b1_S1009 = 1010;
  localparam retro_main_b1_S1010 = 1011;
  localparam retro_main_b1_S1011 = 1012;
  localparam retro_main_b1_S1012 = 1013;
  localparam retro_main_b1_S1013 = 1014;
  localparam retro_main_b1_S1014 = 1015;
  localparam retro_main_b1_S1015 = 1016;
  localparam retro_main_b1_S1016 = 1017;
  localparam retro_main_b1_S1017 = 1018;
  localparam retro_main_b1_S1018 = 1019;
  localparam retro_main_b1_S1019 = 1020;
  localparam retro_main_b1_S1020 = 1021;
  localparam retro_main_b1_S1021 = 1022;
  localparam retro_main_b1_S1022 = 1023;
  localparam retro_main_b1_S1023 = 1024;
  localparam retro_main_b1_S1024 = 1025;
  localparam retro_main_whileexit191_FINISH = 1026;
  localparam retro_main_L1_while2_S0 = 1027;
  localparam retro_main_L1_whilebody3_S0 = 1028;
  localparam retro_main_L1_whilebody3_S1 = 1029;
  localparam retro_main_L1_whilebody3_S2 = 1030;
  localparam retro_main_L1_whilebody3_S3 = 1031;
  localparam retro_main_L1_ifthen9_S0 = 1032;
  localparam retro_main_L1_ifelse177_S0 = 1033;
  localparam retro_main_L1_ifelse177_S1 = 1034;
  localparam retro_main_L1_ifelse177_S2 = 1035;
  localparam retro_main_L1_ifelse177_S3 = 1036;
  localparam retro_main_L1_ifthen16_S0 = 1037;
  localparam retro_main_L1_ifthen20_S0 = 1038;
  localparam retro_main_L1_ifthen20_S1 = 1039;
  localparam retro_main_L1_ifthen24_S0 = 1040;
  localparam retro_main_L1_ifthen24_S1 = 1041;
  localparam retro_main_L1_ifthen24_S2 = 1042;
  localparam retro_main_L1_ifthen24_S3 = 1043;
  localparam retro_main_L1_ifthen28_S0 = 1044;
  localparam retro_main_L1_ifthen32_S0 = 1045;
  localparam retro_main_L1_ifthen32_S1 = 1046;
  localparam retro_main_L1_ifthen32_S2 = 1047;
  localparam retro_main_L1_ifthen32_S3 = 1048;
  localparam retro_main_L1_ifthen36_S0 = 1049;
  localparam retro_main_L1_ifthen36_S1 = 1050;
  localparam retro_main_L1_ifthen36_S2 = 1051;
  localparam retro_main_L1_ifthen36_S3 = 1052;
  localparam retro_main_L1_ifthen40_S0 = 1053;
  localparam retro_main_L1_ifthen44_S0 = 1054;
  localparam retro_main_L1_ifthen44_S1 = 1055;
  localparam retro_main_L1_ifthen48_S0 = 1056;
  localparam retro_main_L1_ifthen48_S1 = 1057;
  localparam retro_main_L1_ifthen48_S2 = 1058;
  localparam retro_main_L1_ifthen48_S3 = 1059;
  localparam retro_main_L1_ifthen48_S4 = 1060;
  localparam retro_main_L1_ifthen52_S0 = 1061;
  localparam retro_main_L1_ifthen56_S0 = 1062;
  localparam retro_main_L1_ifthen60_S0 = 1063;
  localparam retro_main_L1_ifthen64_S0 = 1064;
  localparam retro_main_L1_ifthen68_S0 = 1065;
  localparam retro_main_L1_ifthen72_S0 = 1066;
  localparam retro_main_L1_ifthen81_S0 = 1067;
  localparam retro_main_L1_ifthen81_S1 = 1068;
  localparam retro_main_L1_ifthen81_S2 = 1069;
  localparam retro_main_L1_ifthen81_S3 = 1070;
  localparam retro_main_L1_ifthen81_S4 = 1071;
  localparam retro_main_L1_ifthen85_S0 = 1072;
  localparam retro_main_L1_ifthen85_S1 = 1073;
  localparam retro_main_L1_ifthen85_S2 = 1074;
  localparam retro_main_L1_ifthen85_S3 = 1075;
  localparam retro_main_L1_ifthen85_S4 = 1076;
  localparam retro_main_L1_ifthen89_S0 = 1077;
  localparam retro_main_L1_ifthen89_S1 = 1078;
  localparam retro_main_L1_ifthen89_S2 = 1079;
  localparam retro_main_L1_ifthen89_S3 = 1080;
  localparam retro_main_L1_ifthen89_S4 = 1081;
  localparam retro_main_L1_ifthen93_S0 = 1082;
  localparam retro_main_L1_ifthen93_S2 = 1083;
  localparam retro_main_L1_ifthen97_S0 = 1084;
  localparam retro_main_L1_ifthen97_S2 = 1085;
  localparam retro_main_L1_ifthen97_S3 = 1086;
  localparam retro_main_L1_ifthen97_S4 = 1087;
  localparam retro_main_L1_ifthen97_S5 = 1088;
  localparam retro_main_L1_ifthen101_S0 = 1089;
  localparam retro_main_L1_ifthen101_S2 = 1090;
  localparam retro_main_L1_ifthen101_S3 = 1091;
  localparam retro_main_L1_ifthen101_S4 = 1092;
  localparam retro_main_L1_ifthen101_S5 = 1093;
  localparam retro_main_L1_ifthen105_S0 = 1094;
  localparam retro_main_L1_ifthen105_S2 = 1095;
  localparam retro_main_L1_ifthen105_S3 = 1096;
  localparam retro_main_L1_ifthen105_S4 = 1097;
  localparam retro_main_L1_ifthen105_S5 = 1098;
  localparam retro_main_L1_ifthen109_S0 = 1099;
  localparam retro_main_L1_ifthen109_S2 = 1100;
  localparam retro_main_L1_ifthen109_S3 = 1101;
  localparam retro_main_L1_ifthen109_S4 = 1102;
  localparam retro_main_L1_ifthen109_S5 = 1103;
  localparam retro_main_L1_ifthen113_S0 = 1104;
  localparam retro_main_L1_ifthen113_S2 = 1105;
  localparam retro_main_L1_ifthen113_S3 = 1106;
  localparam retro_main_L1_ifthen113_S4 = 1107;
  localparam retro_main_L1_ifthen113_S5 = 1108;
  localparam retro_main_L1_ifthen117_S0 = 1109;
  localparam retro_main_L1_ifthen121_S0 = 1110;
  localparam retro_main_L1_ifthen125_S0 = 1111;
  localparam retro_main_L1_ifthen125_S3 = 1112;
  localparam retro_main_L1_ifthen129_S0 = 1113;
  localparam retro_main_L1_ifthen129_S1 = 1114;
  localparam retro_main_L1_ifthen133_S0 = 1115;
  localparam retro_main_L1_ifthen133_S3 = 1116;
  localparam retro_main_L1_ifthen133_S4 = 1117;
  localparam retro_main_L1_ifthen133_S5 = 1118;
  localparam retro_main_L1_ifthen133_S6 = 1119;
  localparam retro_main_L1_ifthen133_S7 = 1120;
  localparam retro_main_L1_ifthen137_S0 = 1121;
  localparam retro_main_L1_ifthen137_S1 = 1122;
  localparam retro_main_L1_ifthen218_S0 = 1123;
  localparam retro_main_L1_ifthen220_S0 = 1124;
  localparam retro_main_L1_ifelse221_S0 = 1125;
  localparam retro_main_L1_ifelse221_S3 = 1126;
  localparam retro_main_L1_ifelse221_S4 = 1127;
  localparam retro_main_L1_ifthen304_S0 = 1128;
  localparam retro_main_L1_ifthen304_S3 = 1129;
  localparam retro_main_L1_ifthen316_S0 = 1130;
  localparam retro_main_L1_ifthen317_S0 = 1131;
  localparam retro_main_L1_ifthen317_S7 = 1132;
  localparam retro_main_L1_ifelse318_S0 = 1133;
  localparam retro_main_L1_ifelse318_S1 = 1134;
  localparam retro_main_L1_ifelse325_S0 = 1135;
  localparam retro_main_L1_ifelse325_S1 = 1136;
  localparam retro_main_L1_ifthen328_S0 = 1137;
  localparam retro_main_L1_ifthen328_S1 = 1138;
  localparam retro_main_L1_ifthen328_S3 = 1139;
  localparam retro_main_L1_ifthen328_S4 = 1140;
  localparam retro_main_L1_ifthen328_S5 = 1141;
  localparam retro_main_L1_ifthen328_S6 = 1142;
  localparam retro_main_L1_ifthen334_S0 = 1143;
  localparam retro_main_L1_ifthen334_S4 = 1144;
  localparam retro_main_L1_ifthen334_S5 = 1145;
  localparam retro_main_L1_ifthen334_S6 = 1146;
  localparam retro_main_L1_ifthen334_S7 = 1147;
  localparam retro_main_L1_ifthen341_S0 = 1148;
  localparam retro_main_L1_ifthen341_S7 = 1149;
  localparam retro_main_L1_ifelse342_S0 = 1150;
  localparam retro_main_L1_ifelse342_S1 = 1151;
  localparam retro_main_L1_ifthen345_S0 = 1152;
  localparam retro_main_L1_ifthen345_S1 = 1153;
  localparam retro_main_L1_ifthen345_S4 = 1154;
  localparam retro_main_L1_ifthen345_S5 = 1155;
  localparam retro_main_L1_ifthen345_S6 = 1156;
  localparam retro_main_L1_ifthen345_S7 = 1157;
  localparam retro_main_L1_ifthen351_S0 = 1158;
  localparam retro_main_L1_ifthen351_S4 = 1159;
  localparam retro_main_L1_ifthen351_S5 = 1160;
  localparam retro_main_L1_ifthen351_S6 = 1161;
  localparam retro_main_L1_ifthen351_S7 = 1162;
  localparam retro_main_L1_ifthen358_S0 = 1163;
  localparam retro_main_L1_ifthen358_S7 = 1164;
  localparam retro_main_L1_ifelse359_S0 = 1165;
  localparam retro_main_L1_ifelse359_S1 = 1166;
  localparam retro_main_L1_ifthen362_S0 = 1167;
  localparam retro_main_L1_ifthen362_S1 = 1168;
  localparam retro_main_L1_ifthen362_S4 = 1169;
  localparam retro_main_L1_ifthen362_S5 = 1170;
  localparam retro_main_L1_ifthen362_S6 = 1171;
  localparam retro_main_L1_ifthen362_S7 = 1172;
  localparam retro_main_L1_ifthen368_S0 = 1173;
  localparam retro_main_L1_ifthen368_S4 = 1174;
  localparam retro_main_L1_ifthen368_S5 = 1175;
  localparam retro_main_L1_ifthen368_S6 = 1176;
  localparam retro_main_L1_ifthen368_S7 = 1177;
  localparam retro_main_L1_ifthen375_S0 = 1178;
  localparam retro_main_L1_ifthen375_S7 = 1179;
  localparam retro_main_L1_ifelse376_S0 = 1180;
  localparam retro_main_L1_ifelse376_S1 = 1181;
  localparam retro_main_L1_ifthen379_S0 = 1182;
  localparam retro_main_L1_ifthen379_S1 = 1183;
  localparam retro_main_L1_ifthen379_S5 = 1184;
  localparam retro_main_L1_ifthen379_S6 = 1185;
  localparam retro_main_L1_ifthen379_S7 = 1186;
  localparam retro_main_L1_ifthen379_S8 = 1187;
  localparam retro_main_L1_ifthen385_S0 = 1188;
  localparam retro_main_L1_ifthen385_S5 = 1189;
  localparam retro_main_L1_ifthen385_S6 = 1190;
  localparam retro_main_L1_ifthen385_S7 = 1191;
  localparam retro_main_L1_ifthen385_S8 = 1192;
  localparam retro_main_L1_ifthen392_S0 = 1193;
  localparam retro_main_L1_ifthen392_S7 = 1194;
  localparam retro_main_L1_ifelse393_S0 = 1195;
  localparam retro_main_L1_ifelse393_S1 = 1196;
  localparam retro_main_L1_ifthen396_S0 = 1197;
  localparam retro_main_L1_ifthen398_S0 = 1198;
  localparam retro_main_L1_ifthen399_S0 = 1199;
  localparam retro_main_L1_ifelse404_S0 = 1200;
  localparam retro_main_L1_ifelse404_S1 = 1201;
  localparam retro_main_L1_ifthen407_S0 = 1202;
  localparam retro_main_L1_ifthen407_S5 = 1203;
  localparam retro_main_L1_ifthen407_S6 = 1204;
  localparam retro_main_L1_ifthen407_S7 = 1205;
  localparam retro_main_L1_ifthen407_S8 = 1206;
  localparam retro_main_L1_ifelse413_S0 = 1207;
  localparam retro_main_L1_ifelse413_S5 = 1208;
  localparam retro_main_L1_ifelse413_S6 = 1209;
  localparam retro_main_L1_ifelse413_S7 = 1210;
  localparam retro_main_L1_ifelse413_S8 = 1211;
  localparam retro_main_L1_ifthen478_S0 = 1212;
  localparam retro_main_L1_ifelse490_S0 = 1213;
  localparam retro_main_L1_ifelse490_S1 = 1214;
  localparam retro_main_L1_ifthen140_S0 = 1215;
  localparam retro_main_L1_ifthen140_S1 = 1216;
  localparam retro_main_L1_exit219_S0 = 1217;
  localparam retro_main_L1_ifthen309_S0 = 1218;
  localparam retro_main_L1_ifelse311_S0 = 1219;
  localparam retro_main_L1_ifelse311_S5 = 1220;
  localparam retro_main_L1_ifelse311_S6 = 1221;
  localparam retro_main_L1_ifelse311_S7 = 1222;
  localparam retro_main_L1_ifelse311_S8 = 1223;
  localparam retro_main_L1_exit322_S0 = 1224;
  localparam retro_main_L1_b564_S0 = 1225;
  localparam retro_main_L1_b565_S0 = 1226;
  localparam retro_main_L1_b566_S0 = 1227;
  localparam retro_main_L1_b567_S0 = 1228;
  localparam retro_main_L1_exit397_S0 = 1229;
  localparam retro_main_L1_exit412_S0 = 1230;
  localparam retro_main_L1_ifthen479_S0 = 1231;
  localparam retro_main_L1_ifthen479_S6 = 1232;
  localparam retro_main_L1_ifthen479_S7 = 1233;
  localparam retro_main_L1_ifthen479_S8 = 1234;
  localparam retro_main_L1_ifthen479_S9 = 1235;
  localparam retro_main_L1_ifelse489_S0 = 1236;
  localparam retro_main_L1_ifthen493_S0 = 1237;
  localparam retro_main_L1_ifthen493_S1 = 1238;
  localparam retro_main_L1_ifthen493_S2 = 1239;
  localparam retro_main_L1_ifthen493_S3 = 1240;
  localparam retro_main_L1_exit310_S0 = 1241;
  localparam retro_main_L1_exit310_S1 = 1242;
  localparam retro_main_L1_exit333_S0 = 1243;
  localparam retro_main_L1_exit350_S0 = 1244;
  localparam retro_main_L1_exit367_S0 = 1245;
  localparam retro_main_L1_exit384_S0 = 1246;
  localparam retro_main_L1_b568_S0 = 1247;
  localparam retro_main_L1_exit488_S0 = 1248;
  localparam retro_main_L1_ifthen496_S0 = 1249;
  localparam retro_main_L1_ifthen496_S1 = 1250;
  localparam retro_main_L1_b497_S0 = 1251;
  localparam retro_main_L1_b497_S1 = 1252;
  localparam retro_main_L1_ifthen498_S0 = 1253;
  localparam retro_main_L1_ifthen499_S0 = 1254;
  localparam retro_main_L1_ifelse558_S0 = 1255;
  localparam retro_main_L1_ifelse558_S6 = 1256;
  localparam retro_main_L1_ifelse558_S7 = 1257;
  localparam retro_main_L1_ifelse558_S8 = 1258;
  localparam retro_main_L1_ifelse558_S9 = 1259;
  localparam retro_main_L1_ifthen500_S0 = 1260;
  localparam retro_main_L1_ifthen500_S6 = 1261;
  localparam retro_main_L1_ifthen500_S7 = 1262;
  localparam retro_main_L1_ifthen500_S8 = 1263;
  localparam retro_main_L1_ifthen500_S9 = 1264;
  localparam retro_main_L1_ifthen500_S10 = 1265;
  localparam retro_main_L1_ifthen500_S11 = 1266;
  localparam retro_main_L1_ifthen500_S12 = 1267;
  localparam retro_main_L1_ifelse551_S0 = 1268;
  localparam retro_main_L1_ifelse551_S6 = 1269;
  localparam retro_main_L1_ifelse551_S7 = 1270;
  localparam retro_main_L1_ifelse551_S8 = 1271;
  localparam retro_main_L1_ifelse551_S9 = 1272;
  localparam retro_main_L1_ifelse551_S10 = 1273;
  localparam retro_main_L1_b511_S0 = 1274;
  localparam retro_main_L1_b511_S1 = 1275;
  localparam retro_main_L1_b514_S0 = 1276;
  localparam retro_main_L1_b514_S1 = 1277;
  localparam retro_main_L1_ifthen515_S0 = 1278;
  localparam retro_main_L1_ifthen515_S1 = 1279;
  localparam retro_main_L1_b516_S0 = 1280;
  localparam retro_main_L1_b516_S1 = 1281;
  localparam retro_main_L1_ifthen517_S0 = 1282;
  localparam retro_main_L1_ifthen517_S1 = 1283;
  localparam retro_main_L1_b518_S0 = 1284;
  localparam retro_main_L1_b518_S1 = 1285;
  localparam retro_main_L1_ifthen519_S0 = 1286;
  localparam retro_main_L1_ifthen519_S1 = 1287;
  localparam retro_main_L1_ifthen545_S0 = 1288;
  localparam retro_main_L1_ifthen545_S1 = 1289;
  localparam retro_main_L1_ifthen546_S0 = 1290;
  localparam retro_main_L1_ifthen546_S1 = 1291;
  localparam retro_main_L1_ifthen547_S0 = 1292;
  localparam retro_main_L1_ifthen547_S1 = 1293;
  localparam retro_main_L1_ifthen548_S0 = 1294;
  localparam retro_main_L1_ifthen548_S1 = 1295;
  localparam retro_main_L1_ifthen549_S0 = 1296;
  localparam retro_main_L1_ifthen549_S1 = 1297;
  localparam retro_main_L1_ifthen550_S0 = 1298;
  localparam retro_main_L1_ifthen550_S1 = 1299;
  localparam retro_main_L1_b520_S0 = 1300;
  localparam retro_main_L1_b520_S1 = 1301;
  localparam retro_main_L1_ifthen521_S0 = 1302;
  localparam retro_main_L1_ifthen521_S1 = 1303;
  localparam retro_main_L1_b522_S0 = 1304;
  localparam retro_main_L1_b522_S1 = 1305;
  localparam retro_main_L1_ifthen523_S0 = 1306;
  localparam retro_main_L1_ifthen523_S1 = 1307;
  localparam retro_main_L1_ifthen527_S0 = 1308;
  localparam retro_main_L1_ifthen527_S1 = 1309;
  localparam retro_main_L1_ifthen528_S0 = 1310;
  localparam retro_main_L1_ifthen528_S1 = 1311;
  localparam retro_main_L1_ifthen529_S0 = 1312;
  localparam retro_main_L1_ifthen529_S1 = 1313;
  localparam retro_main_L1_ifthen530_S0 = 1314;
  localparam retro_main_L1_ifthen530_S1 = 1315;
  localparam retro_main_L1_ifthen533_S0 = 1316;
  localparam retro_main_L1_ifthen533_S1 = 1317;
  localparam retro_main_L1_ifthen536_S0 = 1318;
  localparam retro_main_L1_ifthen536_S1 = 1319;
  localparam retro_main_L1_ifthen537_S0 = 1320;
  localparam retro_main_L1_ifthen537_S1 = 1321;
  localparam retro_main_L1_ifthen538_S0 = 1322;
  localparam retro_main_L1_ifthen538_S1 = 1323;
  localparam retro_main_L1_ifthen539_S0 = 1324;
  localparam retro_main_L1_ifthen539_S1 = 1325;
  localparam retro_main_L1_ifthen540_S0 = 1326;
  localparam retro_main_L1_ifthen540_S1 = 1327;
  localparam retro_main_L1_ifthen541_S0 = 1328;
  localparam retro_main_L1_ifthen541_S1 = 1329;
  localparam retro_main_L1_ifthen542_S0 = 1330;
  localparam retro_main_L1_ifthen542_S1 = 1331;
  localparam retro_main_L1_ifthen543_S0 = 1332;
  localparam retro_main_L1_ifthen543_S1 = 1333;
  localparam retro_main_L1_ifthen544_S0 = 1334;
  localparam retro_main_L1_ifthen544_S1 = 1335;
  localparam retro_main_L1_b524_S0 = 1336;
  localparam retro_main_L1_b524_S1 = 1337;
  localparam retro_main_L1_ifthen525_S0 = 1338;
  localparam retro_main_L1_ifthen525_S1 = 1339;
  localparam retro_main_L1_b526_S0 = 1340;
  localparam retro_main_L1_b178_S0 = 1341;
  localparam retro_main_L1_b178_S1 = 1342;
  localparam retro_main_L1_ifthen179_S0 = 1343;
  localparam retro_main_L1_ifthen179_S1 = 1344;
  localparam retro_main_L1_b183_S0 = 1345;
  localparam retro_main_L1_b183_S1 = 1346;
  localparam retro_main_L1_b183_S2 = 1347;
  
  //signals: 
  reg        [31:0] array1007_inl52 [0:1];
  reg        [31:0] array1010 [0:11];
  wire c1000_inl52;
  wire c1001_inl52;
  wire c1002_inl52;
  wire c1003_inl52;
  wire c1004_inl52;
  wire c1005_inl1_inl52;
  wire c1005_inl2_inl52;
  wire c1018_inl39;
  wire c1019_inl39;
  wire c1020_inl39;
  wire c1021_inl38;
  wire c1022_inl38;
  wire c1023_inl38;
  wire c1024_inl37;
  wire c1025_inl37;
  wire c1026_inl37;
  wire c1027_inl36;
  wire c1028_inl36;
  wire c1029_inl36;
  wire c1030_inl35;
  wire c1031_inl35;
  wire c1032_inl35;
  wire c1033_inl33;
  wire c1034_inl33;
  wire c1035_inl33;
  wire c1036_inl13;
  wire c1037_inl13;
  wire c1038_inl34;
  wire c1039_inl34;
  wire c1040_inl34;
  wire c1041;
  wire c1042;
  wire c1043;
  wire c1044;
  wire c1045;
  wire c1046;
  wire c1047;
  wire c1048;
  wire c1049;
  wire c1050;
  wire c1051;
  wire c1052;
  wire c1053;
  wire c1054;
  wire c1055;
  wire c1056;
  wire c1057;
  wire c1058;
  wire c1059;
  wire c1060;
  wire c1061;
  wire c1062;
  wire c1063;
  wire c1064;
  wire c1065;
  wire c1066;
  wire c1067;
  wire c1068;
  wire c1069;
  wire c1070;
  wire c1071;
  wire c1072_inl55;
  wire c1073_inl55;
  wire c1074_inl55;
  wire c1075_inl55;
  wire c1076_inl55;
  wire c1077_inl55;
  wire c1078_inl55;
  wire c1079_inl55;
  wire c1080_inl55;
  wire c1081_inl55;
  wire c1082_inl55;
  wire c1083_inl55;
  wire c1084_inl55;
  wire c1085_inl55;
  wire c1086_inl55;
  wire c1087_inl55;
  wire c1088_inl55;
  wire c1089_inl55;
  wire c1090_inl55;
  wire c1091_inl55;
  wire c1092_inl55;
  wire c1093_inl55;
  wire c1094_inl52;
  wire c1095_inl52;
  wire c1096_inl52;
  wire c1970;
  wire c1971;
  wire c1972;
  wire c1973;
  wire c1974;
  wire c1975;
  wire c1976;
  wire c1977;
  wire c1978;
  wire c1979;
  wire c1980;
  wire c1981;
  wire c1982;
  wire c1983;
  wire c1984;
  wire c1985;
  wire c1986;
  wire c1987;
  wire c1988;
  wire c1989;
  wire c1990;
  wire c1991;
  wire c1992;
  wire c1993;
  wire c1994;
  wire c1995;
  wire c1996;
  wire c1997;
  wire c1998;
  wire c1999;
  wire c2000;
  wire c2001;
  wire c2002;
  wire c2004;
  wire c2005;
  wire c2006;
  wire c2012;
  wire c2013;
  wire c2014;
  wire c2015;
  wire c2016;
  wire c2017;
  wire c2018;
  wire c2019;
  wire c2021;
  wire c2022;
  wire c2023;
  wire c2024;
  wire c2025;
  wire c2026;
  wire c2027;
  wire c2028;
  wire c2029;
  wire c2030;
  wire c2031;
  wire c2032;
  wire c2033;
  wire c2034;
  wire c2035;
  wire c2036;
  wire c2037;
  wire c2038;
  wire c2039;
  wire c2040;
  wire c2041;
  wire c2042;
  wire c2046;
  wire c2047;
  wire c2048;
  wire c2054;
  wire c2055;
  wire c2060;
  wire c2090;
  wire c2091;
  wire c2093;
  wire c2120;
  wire c2124;
  wire c2125;
  wire c2126;
  wire c2127;
  wire c2128;
  wire c2129;
  wire c2130;
  wire c2131;
  wire c2132;
  wire c2133;
  wire c2139;
  wire c2140;
  wire c2146;
  wire c2148;
  wire c2151;
  wire c2152;
  wire c2155;
  wire c2156;
  wire c2166;
  wire c2167;
  wire c2168;
  wire c2169;
  wire c2170;
  wire c2171;
  wire c2172;
  wire c2173;
  wire c2174;
  wire c2175;
  wire c2176;
  wire c2177;
  wire c2178;
  wire c2179;
  wire c2180;
  wire c2181;
  wire c2182;
  wire c2183;
  wire c2184;
  wire c2185;
  wire c2186;
  wire c2187;
  wire c2188;
  wire c2189;
  wire c2190;
  wire c2191;
  wire c2192;
  wire c2193;
  wire c2194;
  wire c2195;
  wire c2196;
  wire c2197;
  wire c2198;
  wire c2199;
  wire c2200;
  wire c2201;
  wire c3337;
  wire c3338;
  wire c3339;
  wire c3340;
  wire c3341;
  wire c3342;
  wire c3343;
  wire c3344;
  wire c3345;
  wire c3346;
  wire c3347;
  wire c3348;
  wire c3349;
  wire c3350;
  wire c3351;
  wire c3352;
  wire c3353;
  wire c3354;
  wire c3355;
  wire c3356;
  wire c3357;
  wire c3358;
  wire c3359;
  wire c3360;
  wire c3361;
  wire c3362;
  wire c3363;
  wire c3364;
  wire c3365;
  wire c3366;
  wire c3367;
  wire c3368;
  wire c3369;
  wire c3370;
  wire c3371;
  wire c3372;
  wire c3373;
  wire c3374;
  wire c3375;
  wire c3376;
  wire c3377;
  wire c3378;
  wire c3379;
  wire c3380;
  wire c3381;
  wire c3382;
  wire c3383;
  wire c3384;
  wire c3385;
  wire c3386;
  wire c3387;
  wire c3388;
  wire c3389;
  wire c3390;
  wire c3391;
  wire c3392;
  wire c3393;
  wire c3394;
  wire c3395;
  wire c3396;
  wire c3397;
  wire c3398;
  wire c3399;
  wire c3400;
  wire c3401;
  wire c3402;
  wire c3403;
  wire c3404;
  wire c3405;
  wire c3406;
  wire c3407;
  wire c3408;
  wire c3409;
  wire c3410;
  wire c3411;
  wire c3412;
  wire c3413;
  wire c3414;
  wire c3415;
  wire c3416;
  wire c3417;
  wire c3418;
  wire c3419;
  wire c3420;
  wire c3421;
  wire c3422;
  wire c3423;
  wire c3424;
  wire c3425;
  wire c3426;
  wire c3427;
  wire c3428;
  wire c3429;
  wire c3430;
  wire c3431;
  wire c3432;
  wire c3433;
  wire c3434;
  wire c3435;
  wire c3436;
  wire c3437;
  wire c3438;
  wire c3439;
  wire c3440;
  wire c3441;
  wire c3442;
  wire c3443;
  wire c3444;
  wire c3445;
  wire c3446;
  wire c3447;
  wire c3448;
  wire c3449;
  wire c3450;
  wire c843_inl40;
  wire c845_inl54;
  wire c846_inl54;
  wire c848_inl39;
  wire c849_inl39;
  wire c850_inl39;
  wire c852_inl38;
  wire c853_inl38;
  wire c854_inl38;
  wire c855_inl38;
  wire c857_inl37;
  wire c858_inl37;
  wire c859_inl37;
  wire c860_inl37;
  wire c862_inl36;
  wire c863_inl36;
  wire c864_inl36;
  wire c865_inl36;
  wire c867_inl35;
  wire c868_inl35;
  wire c869_inl35;
  wire c870_inl35;
  wire c872_inl33;
  wire c873_inl33;
  wire c874_inl33;
  wire c875_inl33;
  wire c876_inl33;
  wire c877_inl33;
  wire c879_inl13;
  wire c880_inl13;
  wire c882_inl34;
  wire c883_inl34;
  wire c884_inl34;
  wire c886;
  wire c887;
  wire c888;
  wire c889;
  wire c890;
  wire c891;
  wire c892;
  wire c893;
  wire c894;
  wire c895;
  wire c896;
  wire c897;
  wire c898;
  wire c899;
  wire c900;
  wire c901;
  wire c902;
  wire c903;
  wire c904;
  wire c905;
  wire c906;
  wire c907;
  wire c908;
  wire c909;
  wire c910;
  wire c911;
  wire c912;
  wire c913;
  wire c914;
  wire c915;
  wire c916;
  wire c917;
  wire c918;
  wire c919;
  wire c920;
  wire c921;
  wire c924;
  wire c927;
  wire c930_inl55;
  wire c933_inl55;
  wire c935_inl55;
  wire c936_inl55;
  wire c937_inl55;
  wire c938_inl55;
  wire c939_inl55;
  wire c942_inl55;
  wire c944_inl55;
  wire c946_inl55;
  wire c948_inl55;
  wire c950_inl55;
  wire c952_inl55;
  wire c954_inl55;
  wire c956_inl55;
  wire c958_inl55;
  wire c960_inl55;
  wire c962_inl55;
  wire c964_inl55;
  wire c966_inl55;
  wire c968_inl55;
  wire c970_inl55;
  wire c972_inl55;
  wire c974_inl55;
  wire c976_inl55;
  wire c978_inl55;
  wire c980_inl55;
  wire c982_inl55;
  wire c984_inl55;
  wire c986_inl55;
  wire c988_inl55;
  wire c990_inl55;
  wire c992_inl55;
  wire c996_inl52;
  wire c997_inl52;
  wire c998_inl52;
  wire c999_inl52;
  wire done_flag13;
  wire exec_result135;
  wire exec_result346;
  wire exec_result357;
  wire exec_result367;
  wire exec_result377;
  wire exec_result387;
  wire exec_result396;
  wire exec_result404;
  wire exec_result545;
  wire        [31:0] retro_divmod_result522 [0:1];
  wire t2771;
  wire t2778;
  wire t2785;
  wire t2792;
  wire t2829;
  wire wr_flag4;
  wire wr_flag6;
  reg done_flag2;
  reg exec_result336;
  reg        [10:0] retro_main_state;
  reg wr_flag2;
  wire signed [31:0] address0_pos3;
  wire signed [31:0] address0_pos4;
  wire signed [31:0] address0_pos5;
  wire signed [31:0] address0_pos6;
  wire signed [31:0] address0_pos7;
  wire signed [31:0] address0_pos8;
  wire signed [31:0] address0_pos9;
  wire signed [31:0] address0_second7;
  wire signed [31:0] address0_second9;
  wire signed [31:0] address0_top7;
  wire signed [31:0] address0_top9;
  wire signed [31:0] ip15;
  wire signed [31:0] ip16;
  wire signed [31:0] ip17;
  wire signed [31:0] ip18;
  wire signed [31:0] ip_inl554;
  wire signed [31:0] jump0_ip3;
  wire signed [31:0] jump0_ip4;
  wire signed [31:0] jump0_ip5;
  wire signed [31:0] jump0_ip6;
  wire signed [31:0] jump0_phase7;
  wire signed [31:0] jump0_phase8;
  wire signed [31:0] jump_eq0_a4;
  wire signed [31:0] jump_eq0_a5;
  wire signed [31:0] jump_eq0_ip3;
  wire signed [31:0] jump_eq0_ip4;
  wire signed [31:0] jump_eq0_ip5;
  wire signed [31:0] jump_eq0_ip6;
  wire signed [31:0] jump_eq0_phase8;
  wire signed [31:0] jump_eq0_phase9;
  wire signed [31:0] jump_ge0_a4;
  wire signed [31:0] jump_ge0_a5;
  wire signed [31:0] jump_ge0_ip3;
  wire signed [31:0] jump_ge0_ip4;
  wire signed [31:0] jump_ge0_ip5;
  wire signed [31:0] jump_ge0_ip6;
  wire signed [31:0] jump_ge0_phase8;
  wire signed [31:0] jump_ge0_phase9;
  wire signed [31:0] jump_le0_a4;
  wire signed [31:0] jump_le0_a5;
  wire signed [31:0] jump_le0_ip3;
  wire signed [31:0] jump_le0_ip4;
  wire signed [31:0] jump_le0_ip5;
  wire signed [31:0] jump_le0_ip6;
  wire signed [31:0] jump_le0_phase8;
  wire signed [31:0] jump_le0_phase9;
  wire signed [31:0] jump_ne0_a4;
  wire signed [31:0] jump_ne0_a5;
  wire signed [31:0] jump_ne0_ip3;
  wire signed [31:0] jump_ne0_ip4;
  wire signed [31:0] jump_ne0_ip5;
  wire signed [31:0] jump_ne0_ip6;
  wire signed [31:0] jump_ne0_phase8;
  wire signed [31:0] jump_ne0_phase9;
  wire signed [31:0] lit0_ip3;
  wire signed [31:0] lit0_ip4;
  wire signed [31:0] lit0_ip5;
  wire signed [31:0] lit0_phase6;
  wire signed [31:0] lit0_phase7;
  wire signed [31:0] loop0_ip3;
  wire signed [31:0] loop0_ip4;
  wire signed [31:0] loop0_ip5;
  wire signed [31:0] loop0_ip6;
  wire signed [31:0] loop0_phase8;
  wire signed [31:0] loop0_phase9;
  wire signed [31:0] opcode4;
  wire signed [31:0] point0_ip5;
  wire signed [31:0] point0_ip6;
  wire signed [31:0] point0_ip_saved4;
  wire signed [31:0] point0_ip_saved5;
  wire signed [31:0] point0_phase7;
  wire signed [31:0] point0_phase8;
  wire signed [31:0] q_inl522;
  wire signed [31:0] q_inl523;
  wire signed [31:0] q_inl524;
  wire signed [31:0] q_inl525;
  wire signed [31:0] r_inl522;
  wire signed [31:0] r_inl523;
  wire signed [31:0] r_inl524;
  wire signed [31:0] r_inl525;
  wire signed [31:0] stack0_pos10;
  wire signed [31:0] stack0_pos11;
  wire signed [31:0] stack0_pos12;
  wire signed [31:0] stack0_pos13;
  wire signed [31:0] stack0_pos14;
  wire signed [31:0] stack0_pos15;
  wire signed [31:0] stack0_pos16;
  wire signed [31:0] stack0_pos17;
  wire signed [31:0] stack0_pos18;
  wire signed [31:0] stack0_pos19;
  wire signed [31:0] stack0_pos20;
  wire signed [31:0] stack0_pos21;
  wire signed [31:0] stack0_pos22;
  wire signed [31:0] stack0_pos23;
  wire signed [31:0] stack0_pos24;
  wire signed [31:0] stack0_pos25;
  wire signed [31:0] stack0_pos26;
  wire signed [31:0] stack0_pos27;
  wire signed [31:0] stack0_pos28;
  wire signed [31:0] stack0_pos29;
  wire signed [31:0] stack0_pos30;
  wire signed [31:0] stack0_pos31;
  wire signed [31:0] stack0_pos32;
  wire signed [31:0] stack0_pos33;
  wire signed [31:0] stack0_pos34;
  wire signed [31:0] stack0_pos35;
  wire signed [31:0] stack0_pos36;
  wire signed [31:0] stack0_pos37;
  wire signed [31:0] stack0_pos38;
  wire signed [31:0] stack0_pos39;
  wire signed [31:0] stack0_pos3;
  wire signed [31:0] stack0_pos40;
  wire signed [31:0] stack0_pos41;
  wire signed [31:0] stack0_pos42;
  wire signed [31:0] stack0_pos43;
  wire signed [31:0] stack0_pos4;
  wire signed [31:0] stack0_pos5;
  wire signed [31:0] stack0_pos6;
  wire signed [31:0] stack0_pos7;
  wire signed [31:0] stack0_pos8;
  wire signed [31:0] stack0_pos9;
  wire signed [31:0] stack0_second11;
  wire signed [31:0] stack0_second14;
  wire signed [31:0] stack0_second17;
  wire signed [31:0] stack0_second20;
  wire signed [31:0] stack0_second23;
  wire signed [31:0] stack0_second26;
  wire signed [31:0] stack0_second30;
  wire signed [31:0] stack0_second37;
  wire signed [31:0] stack0_second43;
  wire signed [31:0] stack0_second44;
  wire signed [31:0] stack0_second45;
  wire signed [31:0] stack0_second4;
  wire signed [31:0] stack0_top10;
  wire signed [31:0] stack0_top12;
  wire signed [31:0] stack0_top15;
  wire signed [31:0] stack0_top18;
  wire signed [31:0] stack0_top21;
  wire signed [31:0] stack0_top24;
  wire signed [31:0] stack0_top26;
  wire signed [31:0] stack0_top31;
  wire signed [31:0] stack0_top33;
  wire signed [31:0] stack0_top35;
  wire signed [31:0] stack0_top36;
  wire signed [31:0] stack0_top38;
  wire signed [31:0] stack0_top40;
  wire signed [31:0] stack0_top42;
  wire signed [31:0] stack0_top44;
  wire signed [31:0] stack0_top46;
  wire signed [31:0] stack0_top48;
  wire signed [31:0] stack0_top49;
  wire signed [31:0] stack0_top4;
  wire signed [31:0] stack0_top50;
  wire signed [31:0] stack0_top58;
  wire signed [31:0] stack0_top59;
  wire signed [31:0] t1006_inl1_inl52;
  wire signed [31:0] t1006_inl2_inl52;
  wire signed [31:0] t2774;
  wire signed [31:0] t2781;
  wire signed [31:0] t2788;
  wire signed [31:0] t2795;
  wire signed [31:0] t2830;
  wire signed [31:0] t2831;
  wire signed [31:0] t839_inl14;
  wire signed [31:0] t839_inl15;
  wire signed [31:0] t839_inl16;
  wire signed [31:0] t839_inl17;
  wire signed [31:0] t839_inl1_inl13;
  wire signed [31:0] t842_inl18;
  wire signed [31:0] t842_inl19;
  wire signed [31:0] t842_inl1_inl35;
  wire signed [31:0] t842_inl1_inl36;
  wire signed [31:0] t842_inl1_inl37;
  wire signed [31:0] t842_inl1_inl38;
  wire signed [31:0] t842_inl1_inl40;
  wire signed [31:0] t842_inl1_inl54;
  wire signed [31:0] t842_inl20;
  wire signed [31:0] t842_inl21;
  wire signed [31:0] t842_inl22;
  wire signed [31:0] t842_inl23;
  wire signed [31:0] t842_inl24;
  wire signed [31:0] t842_inl25;
  wire signed [31:0] t842_inl26;
  wire signed [31:0] t842_inl27;
  wire signed [31:0] t842_inl28;
  wire signed [31:0] t842_inl29;
  wire signed [31:0] t842_inl2_inl33;
  wire signed [31:0] t842_inl2_inl35;
  wire signed [31:0] t842_inl2_inl36;
  wire signed [31:0] t842_inl2_inl37;
  wire signed [31:0] t842_inl2_inl38;
  wire signed [31:0] t842_inl2_inl40;
  wire signed [31:0] t842_inl2_inl54;
  wire signed [31:0] t842_inl2_inl55;
  wire signed [31:0] t842_inl30;
  wire signed [31:0] t842_inl31;
  wire signed [31:0] t842_inl3_inl55;
  wire signed [31:0] t842_inl4_inl55;
  wire signed [31:0] wr_mem_addr4;
  wire signed [31:0] wr_mem_data4;
  wire signed [31:0] write_point0_addr4;
  wire signed [31:0] write_point0_addr5;
  wire signed [31:0] write_point0_data4;
  wire signed [31:0] write_point0_data5;
  wire signed [31:0] write_point0_ip4;
  wire signed [31:0] write_point0_ip5;
  wire signed [31:0] write_point0_phase5;
  wire signed [31:0] write_point0_phase6;
  wire signed [31:0] zero_pop_return0_ip5;
  wire signed [31:0] zero_pop_return0_ip6;
  wire signed [31:0] zero_pop_return0_phase5;
  wire signed [31:0] zero_pop_return0_phase6;
  reg signed [31:0] address0_pos2;
  reg signed [31:0] address0_second2;
  reg signed [31:0] address0_second4;
  reg signed [31:0] address0_second5;
  reg signed [31:0] address0_second6;
  reg signed [31:0] address0_top2;
  reg signed [31:0] ip2;
  reg signed [31:0] jump0_ip2;
  reg signed [31:0] jump0_phase2;
  reg signed [31:0] jump_eq0_a2;
  reg signed [31:0] jump_eq0_ip2;
  reg signed [31:0] jump_eq0_phase2;
  reg signed [31:0] jump_ge0_a2;
  reg signed [31:0] jump_ge0_ip2;
  reg signed [31:0] jump_ge0_phase2;
  reg signed [31:0] jump_le0_a2;
  reg signed [31:0] jump_le0_ip2;
  reg signed [31:0] jump_le0_phase2;
  reg signed [31:0] jump_ne0_a2;
  reg signed [31:0] jump_ne0_ip2;
  reg signed [31:0] jump_ne0_phase2;
  reg signed [31:0] lit0_ip2;
  reg signed [31:0] lit0_phase2;
  reg signed [31:0] loop0_ip2;
  reg signed [31:0] loop0_phase2;
  reg signed [31:0] mem_data;
  reg signed [31:0] opcode2;
  reg signed [31:0] point0_ip2;
  reg signed [31:0] point0_ip_saved2;
  reg signed [31:0] point0_phase2;
  reg signed [31:0] stack0_pos2;
  reg signed [31:0] stack0_second10;
  reg signed [31:0] stack0_second12;
  reg signed [31:0] stack0_second13;
  reg signed [31:0] stack0_second15;
  reg signed [31:0] stack0_second16;
  reg signed [31:0] stack0_second18;
  reg signed [31:0] stack0_second19;
  reg signed [31:0] stack0_second21;
  reg signed [31:0] stack0_second22;
  reg signed [31:0] stack0_second24;
  reg signed [31:0] stack0_second25;
  reg signed [31:0] stack0_second27;
  reg signed [31:0] stack0_second28;
  reg signed [31:0] stack0_second29;
  reg signed [31:0] stack0_second2;
  reg signed [31:0] stack0_second31;
  reg signed [31:0] stack0_second32;
  reg signed [31:0] stack0_second33;
  reg signed [31:0] stack0_second34;
  reg signed [31:0] stack0_second35;
  reg signed [31:0] stack0_second36;
  reg signed [31:0] stack0_second38;
  reg signed [31:0] stack0_second39;
  reg signed [31:0] stack0_second40;
  reg signed [31:0] stack0_second41;
  reg signed [31:0] stack0_second42;
  reg signed [31:0] stack0_second6;
  reg signed [31:0] stack0_second8;
  reg signed [31:0] stack0_top2;
  reg signed [31:0] stack0_top51;
  reg signed [31:0] t11;
  reg signed [31:0] t926;
  reg signed [31:0] t928;
  reg signed [31:0] t929_inl55;
  reg signed [31:0] t932_inl55;
  reg signed [31:0] t934_inl55;
  reg signed [31:0] t941_inl55;
  reg signed [31:0] t943_inl55;
  reg signed [31:0] t945_inl55;
  reg signed [31:0] t947_inl55;
  reg signed [31:0] t949_inl55;
  reg signed [31:0] t951_inl55;
  reg signed [31:0] t953_inl55;
  reg signed [31:0] t955_inl55;
  reg signed [31:0] t957_inl55;
  reg signed [31:0] t959_inl55;
  reg signed [31:0] t961_inl55;
  reg signed [31:0] t963_inl55;
  reg signed [31:0] t965_inl55;
  reg signed [31:0] t967_inl55;
  reg signed [31:0] t969_inl55;
  reg signed [31:0] t971_inl55;
  reg signed [31:0] t973_inl55;
  reg signed [31:0] t975_inl55;
  reg signed [31:0] t977_inl55;
  reg signed [31:0] t979_inl55;
  reg signed [31:0] t981_inl55;
  reg signed [31:0] t983_inl55;
  reg signed [31:0] t985_inl55;
  reg signed [31:0] t987_inl55;
  reg signed [31:0] t989_inl55;
  reg signed [31:0] t991_inl55;
  reg signed [31:0] wr_mem_addr2;
  reg signed [31:0] wr_mem_data2;
  reg signed [31:0] write_point0_addr2;
  reg signed [31:0] write_point0_data2;
  reg signed [31:0] write_point0_ip2;
  reg signed [31:0] write_point0_phase2;
  reg signed [31:0] zero_pop_return0_ip2;
  reg signed [31:0] zero_pop_return0_phase2;
  //signals: _address
  wire        [10:0] _address_len;
  wire        [31:0] _address_q;
  reg        [10:0] _address_addr;
  reg        [31:0] _address_d;
  reg _address_req;
  reg _address_we;
  //signals: _stack
  wire        [7:0] _stack_len;
  wire        [31:0] _stack_q;
  reg        [7:0] _stack_addr;
  reg        [31:0] _stack_d;
  reg _stack_req;
  reg _stack_we;
  //signals: io_ports
  wire        [4:0] io_ports_len;
  wire        [31:0] io_ports_q;
  reg        [4:0] io_ports_addr;
  reg        [31:0] io_ports_d;
  reg io_ports_req;
  reg io_ports_we;
  //signals: memory
  wire        [14:0] memory_len;
  wire        [31:0] memory_q;
  reg        [14:0] memory_addr;
  reg        [31:0] memory_d;
  reg memory_req;
  reg memory_we;
  //signals: ram
  wire        [7:0] array1008_ram_addr;
  wire        [31:0] array1008_ram_d;
  wire        [7:0] array1008_ram_len;
  wire        [31:0] array1008_ram_q;
  wire array1008_ram_we;
  wire        [10:0] array1009_ram_addr;
  wire        [31:0] array1009_ram_d;
  wire        [10:0] array1009_ram_len;
  wire        [31:0] array1009_ram_q;
  wire array1009_ram_we;
  //combinations: 
  assign address0_pos3 = (address0_pos2 + 1);
  assign address0_pos4 = (address0_pos2 - 1);
  assign address0_pos5 = (address0_pos2 - 1);
  assign address0_pos6 = (address0_pos2 - 1);
  assign address0_pos7 = c2090 ? address0_pos6 : c2091 ? address0_pos2 : c2055 ? address0_pos2 : 'bz;
  assign address0_pos8 = (address0_pos2 + 1);
  assign address0_pos9 = (c1971 && c889) ? address0_pos2 : ((c2004 || c2005) || c2006) ? address0_pos2 : c1974 ? address0_pos2 : c1975 ? address0_pos2 : c1976 ? address0_pos2 : c1977 ? address0_pos3 : c1978 ? address0_pos4 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? address0_pos2 : (((c2019 || c2017) || c2018) || c2016) ? address0_pos2 : c1981 ? address0_pos5 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? address0_pos2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? address0_pos2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? address0_pos2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? address0_pos2 : (((c2038 || c2040) || c2037) || c2039) ? address0_pos2 : (c2041 || c2042) ? address0_pos2 : c1988 ? address0_pos2 : c1989 ? address0_pos2 : c1990 ? address0_pos2 : c1991 ? address0_pos2 : c1992 ? address0_pos2 : c1993 ? address0_pos2 : c1994 ? address0_pos2 : c1995 ? address0_pos2 : c1996 ? address0_pos2 : ((c2055 || c2091) || c2090) ? address0_pos7 : c1998 ? address0_pos2 : c1999 ? address0_pos2 : c2000 ? address0_pos2 : c2001 ? address0_pos2 : (c2199 || c2198) ? address0_pos2 : (c2002 && !c927) ? address0_pos2 : c1972 ? address0_pos8 : 'bz;
  assign address0_second7 = c2090 ? address0_second6 : c2091 ? address0_second2 : c2055 ? address0_second2 : 'bz;
  assign address0_second9 = (c1971 && c889) ? address0_second2 : ((c2004 || c2005) || c2006) ? address0_second2 : c1974 ? address0_second2 : c1975 ? address0_second2 : c1976 ? address0_second2 : c1977 ? address0_top2 : c1978 ? address0_second4 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? address0_second2 : (((c2019 || c2017) || c2018) || c2016) ? address0_second2 : c1981 ? address0_second5 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? address0_second2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? address0_second2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? address0_second2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? address0_second2 : (((c2038 || c2040) || c2037) || c2039) ? address0_second2 : (c2041 || c2042) ? address0_second2 : c1988 ? address0_second2 : c1989 ? address0_second2 : c1990 ? address0_second2 : c1991 ? address0_second2 : c1992 ? address0_second2 : c1993 ? address0_second2 : c1994 ? address0_second2 : c1995 ? address0_second2 : c1996 ? address0_second2 : ((c2055 || c2091) || c2090) ? address0_second7 : c1998 ? address0_second2 : c1999 ? address0_second2 : c2000 ? address0_second2 : c2001 ? address0_second2 : (c2199 || c2198) ? address0_second2 : (c2002 && !c927) ? address0_second2 : c1972 ? address0_top2 : 'bz;
  assign address0_top7 = c2090 ? address0_second2 : c2091 ? address0_top2 : c2055 ? address0_top2 : 'bz;
  assign address0_top9 = (c1971 && c889) ? address0_top2 : ((c2004 || c2005) || c2006) ? address0_top2 : c1974 ? address0_top2 : c1975 ? address0_top2 : c1976 ? address0_top2 : c1977 ? stack0_top2 : c1978 ? address0_second2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? address0_top2 : (((c2019 || c2017) || c2018) || c2016) ? address0_top2 : c1981 ? address0_second2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? address0_top2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? address0_top2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? address0_top2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? address0_top2 : (((c2038 || c2040) || c2037) || c2039) ? address0_top2 : (c2041 || c2042) ? address0_top2 : c1988 ? address0_top2 : c1989 ? address0_top2 : c1990 ? address0_top2 : c1991 ? address0_top2 : c1992 ? address0_top2 : c1993 ? address0_top2 : c1994 ? address0_top2 : c1995 ? address0_top2 : c1996 ? address0_top2 : ((c2055 || c2091) || c2090) ? address0_top7 : c1998 ? address0_top2 : c1999 ? address0_top2 : c2000 ? address0_top2 : c2001 ? address0_top2 : (c2199 || c2198) ? address0_top2 : (c2002 && !c927) ? address0_top2 : c1972 ? ip2 : 'bz;
  assign c1000_inl52 = (stack0_top2 < 0);
  assign c1001_inl52 = (c999_inl52 && c1000_inl52);
  assign c1002_inl52 = (stack0_second2 < 0);
  assign c1003_inl52 = (stack0_top2 > 0);
  assign c1004_inl52 = (c1002_inl52 && c1003_inl52);
  assign c1005_inl1_inl52 = (stack0_second2 < 0);
  assign c1005_inl2_inl52 = (stack0_top2 < 0);
  assign c1018_inl39 = (!c848_inl39 && c849_inl39);
  assign c1019_inl39 = ((!c848_inl39 && !c849_inl39) && c850_inl39);
  assign c1020_inl39 = ((!c848_inl39 && !c849_inl39) && !c850_inl39);
  assign c1021_inl38 = (!c852_inl38 && c853_inl38);
  assign c1022_inl38 = ((!c852_inl38 && !c853_inl38) && c854_inl38);
  assign c1023_inl38 = ((!c852_inl38 && !c853_inl38) && !c854_inl38);
  assign c1024_inl37 = (!c857_inl37 && c858_inl37);
  assign c1025_inl37 = ((!c857_inl37 && !c858_inl37) && c859_inl37);
  assign c1026_inl37 = ((!c857_inl37 && !c858_inl37) && !c859_inl37);
  assign c1027_inl36 = (!c862_inl36 && c863_inl36);
  assign c1028_inl36 = ((!c862_inl36 && !c863_inl36) && c864_inl36);
  assign c1029_inl36 = ((!c862_inl36 && !c863_inl36) && !c864_inl36);
  assign c1030_inl35 = (!c867_inl35 && c868_inl35);
  assign c1031_inl35 = ((!c867_inl35 && !c868_inl35) && c869_inl35);
  assign c1032_inl35 = ((!c867_inl35 && !c868_inl35) && !c869_inl35);
  assign c1033_inl33 = (!c872_inl33 && c873_inl33);
  assign c1034_inl33 = ((!c872_inl33 && !c873_inl33) && c874_inl33);
  assign c1035_inl33 = ((!c872_inl33 && !c873_inl33) && !c874_inl33);
  assign c1036_inl13 = (!c879_inl13 && c880_inl13);
  assign c1037_inl13 = (!c879_inl13 && !c880_inl13);
  assign c1038_inl34 = (!c882_inl34 && c883_inl34);
  assign c1039_inl34 = ((!c882_inl34 && !c883_inl34) && c884_inl34);
  assign c1040_inl34 = ((!c882_inl34 && !c883_inl34) && !c884_inl34);
  assign c1041 = (!c889 && c890);
  assign c1042 = ((!c889 && !c890) && c891);
  assign c1043 = (((!c889 && !c890) && !c891) && c892);
  assign c1044 = ((((!c889 && !c890) && !c891) && !c892) && c893);
  assign c1045 = (((((!c889 && !c890) && !c891) && !c892) && !c893) && c894);
  assign c1046 = ((((((!c889 && !c890) && !c891) && !c892) && !c893) && !c894) && c895);
  assign c1047 = (((((((!c889 && !c890) && !c891) && !c892) && !c893) && !c894) && !c895) && c896);
  assign c1048 = ((((((((!c889 && !c890) && !c891) && !c892) && !c893) && !c894) && !c895) && !c896) && c897);
  assign c1049 = (((((((((!c889 && !c890) && !c891) && !c892) && !c893) && !c894) && !c895) && !c896) && !c897) && c898);
  assign c1050 = ((((((((((!c889 && !c890) && !c891) && !c892) && !c893) && !c894) && !c895) && !c896) && !c897) && !c898) && c899);
  assign c1051 = (((((((((((!c889 && !c890) && !c891) && !c892) && !c893) && !c894) && !c895) && !c896) && !c897) && !c898) && !c899) && c900);
  assign c1052 = ((((((((((((!c889 && !c890) && !c891) && !c892) && !c893) && !c894) && !c895) && !c896) && !c897) && !c898) && !c899) && !c900) && c901);
  assign c1053 = (((((((((((((!c889 && !c890) && !c891) && !c892) && !c893) && !c894) && !c895) && !c896) && !c897) && !c898) && !c899) && !c900) && !c901) && c902);
  assign c1054 = ((((((((((((((!c889 && !c890) && !c891) && !c892) && !c893) && !c894) && !c895) && !c896) && !c897) && !c898) && !c899) && !c900) && !c901) && !c902) && c903);
  assign c1055 = (((((((((((((((!c889 && !c890) && !c891) && !c892) && !c893) && !c894) && !c895) && !c896) && !c897) && !c898) && !c899) && !c900) && !c901) && !c902) && !c903) && c904);
  assign c1056 = ((((((((((((((((!c889 && !c890) && !c891) && !c892) && !c893) && !c894) && !c895) && !c896) && !c897) && !c898) && !c899) && !c900) && !c901) && !c902) && !c903) && !c904) && c905);
  assign c1057 = (((((((((((((((((!c889 && !c890) && !c891) && !c892) && !c893) && !c894) && !c895) && !c896) && !c897) && !c898) && !c899) && !c900) && !c901) && !c902) && !c903) && !c904) && !c905) && c906);
  assign c1058 = ((((((((((((((((((!c889 && !c890) && !c891) && !c892) && !c893) && !c894) && !c895) && !c896) && !c897) && !c898) && !c899) && !c900) && !c901) && !c902) && !c903) && !c904) && !c905) && !c906) && c907);
  assign c1059 = (((((((((((((((((((!c889 && !c890) && !c891) && !c892) && !c893) && !c894) && !c895) && !c896) && !c897) && !c898) && !c899) && !c900) && !c901) && !c902) && !c903) && !c904) && !c905) && !c906) && !c907) && c908);
  assign c1060 = ((((((((((((((((((((!c889 && !c890) && !c891) && !c892) && !c893) && !c894) && !c895) && !c896) && !c897) && !c898) && !c899) && !c900) && !c901) && !c902) && !c903) && !c904) && !c905) && !c906) && !c907) && !c908) && c909);
  assign c1061 = (((((((((((((((((((((!c889 && !c890) && !c891) && !c892) && !c893) && !c894) && !c895) && !c896) && !c897) && !c898) && !c899) && !c900) && !c901) && !c902) && !c903) && !c904) && !c905) && !c906) && !c907) && !c908) && !c909) && c910);
  assign c1062 = ((((((((((((((((((((((!c889 && !c890) && !c891) && !c892) && !c893) && !c894) && !c895) && !c896) && !c897) && !c898) && !c899) && !c900) && !c901) && !c902) && !c903) && !c904) && !c905) && !c906) && !c907) && !c908) && !c909) && !c910) && c911);
  assign c1063 = (((((((((((((((((((((((!c889 && !c890) && !c891) && !c892) && !c893) && !c894) && !c895) && !c896) && !c897) && !c898) && !c899) && !c900) && !c901) && !c902) && !c903) && !c904) && !c905) && !c906) && !c907) && !c908) && !c909) && !c910) && !c911) && c912);
  assign c1064 = ((((((((((((((((((((((((!c889 && !c890) && !c891) && !c892) && !c893) && !c894) && !c895) && !c896) && !c897) && !c898) && !c899) && !c900) && !c901) && !c902) && !c903) && !c904) && !c905) && !c906) && !c907) && !c908) && !c909) && !c910) && !c911) && !c912) && c913);
  assign c1065 = (((((((((((((((((((((((((!c889 && !c890) && !c891) && !c892) && !c893) && !c894) && !c895) && !c896) && !c897) && !c898) && !c899) && !c900) && !c901) && !c902) && !c903) && !c904) && !c905) && !c906) && !c907) && !c908) && !c909) && !c910) && !c911) && !c912) && !c913) && c914);
  assign c1066 = ((((((((((((((((((((((((((!c889 && !c890) && !c891) && !c892) && !c893) && !c894) && !c895) && !c896) && !c897) && !c898) && !c899) && !c900) && !c901) && !c902) && !c903) && !c904) && !c905) && !c906) && !c907) && !c908) && !c909) && !c910) && !c911) && !c912) && !c913) && !c914) && c915);
  assign c1067 = (((((((((((((((((((((((((((!c889 && !c890) && !c891) && !c892) && !c893) && !c894) && !c895) && !c896) && !c897) && !c898) && !c899) && !c900) && !c901) && !c902) && !c903) && !c904) && !c905) && !c906) && !c907) && !c908) && !c909) && !c910) && !c911) && !c912) && !c913) && !c914) && !c915) && c916);
  assign c1068 = ((((((((((((((((((((((((((((!c889 && !c890) && !c891) && !c892) && !c893) && !c894) && !c895) && !c896) && !c897) && !c898) && !c899) && !c900) && !c901) && !c902) && !c903) && !c904) && !c905) && !c906) && !c907) && !c908) && !c909) && !c910) && !c911) && !c912) && !c913) && !c914) && !c915) && !c916) && c917);
  assign c1069 = (((((((((((((((((((((((((((((!c889 && !c890) && !c891) && !c892) && !c893) && !c894) && !c895) && !c896) && !c897) && !c898) && !c899) && !c900) && !c901) && !c902) && !c903) && !c904) && !c905) && !c906) && !c907) && !c908) && !c909) && !c910) && !c911) && !c912) && !c913) && !c914) && !c915) && !c916) && !c917) && c918);
  assign c1070 = ((((((((((((((((((((((((((((((!c889 && !c890) && !c891) && !c892) && !c893) && !c894) && !c895) && !c896) && !c897) && !c898) && !c899) && !c900) && !c901) && !c902) && !c903) && !c904) && !c905) && !c906) && !c907) && !c908) && !c909) && !c910) && !c911) && !c912) && !c913) && !c914) && !c915) && !c916) && !c917) && !c918) && c919);
  assign c1071 = ((((((((((((((((((((((((((((((!c889 && !c890) && !c891) && !c892) && !c893) && !c894) && !c895) && !c896) && !c897) && !c898) && !c899) && !c900) && !c901) && !c902) && !c903) && !c904) && !c905) && !c906) && !c907) && !c908) && !c909) && !c910) && !c911) && !c912) && !c913) && !c914) && !c915) && !c916) && !c917) && !c918) && !c919);
  assign c1072_inl55 = (!c946_inl55 && c948_inl55);
  assign c1073_inl55 = ((!c946_inl55 && !c948_inl55) && c950_inl55);
  assign c1074_inl55 = (((!c946_inl55 && !c948_inl55) && !c950_inl55) && c952_inl55);
  assign c1075_inl55 = ((((!c946_inl55 && !c948_inl55) && !c950_inl55) && !c952_inl55) && c954_inl55);
  assign c1076_inl55 = (((((!c946_inl55 && !c948_inl55) && !c950_inl55) && !c952_inl55) && !c954_inl55) && c956_inl55);
  assign c1077_inl55 = ((((((!c946_inl55 && !c948_inl55) && !c950_inl55) && !c952_inl55) && !c954_inl55) && !c956_inl55) && c958_inl55);
  assign c1078_inl55 = ((((((!c946_inl55 && !c948_inl55) && !c950_inl55) && !c952_inl55) && !c954_inl55) && !c956_inl55) && !c958_inl55);
  assign c1079_inl55 = (!c962_inl55 && c964_inl55);
  assign c1080_inl55 = ((!c962_inl55 && !c964_inl55) && c966_inl55);
  assign c1081_inl55 = (((!c962_inl55 && !c964_inl55) && !c966_inl55) && c968_inl55);
  assign c1082_inl55 = ((((!c962_inl55 && !c964_inl55) && !c966_inl55) && !c968_inl55) && c970_inl55);
  assign c1083_inl55 = (((((!c962_inl55 && !c964_inl55) && !c966_inl55) && !c968_inl55) && !c970_inl55) && c972_inl55);
  assign c1084_inl55 = ((((((!c962_inl55 && !c964_inl55) && !c966_inl55) && !c968_inl55) && !c970_inl55) && !c972_inl55) && c974_inl55);
  assign c1085_inl55 = (((((((!c962_inl55 && !c964_inl55) && !c966_inl55) && !c968_inl55) && !c970_inl55) && !c972_inl55) && !c974_inl55) && c976_inl55);
  assign c1086_inl55 = ((((((((!c962_inl55 && !c964_inl55) && !c966_inl55) && !c968_inl55) && !c970_inl55) && !c972_inl55) && !c974_inl55) && !c976_inl55) && c978_inl55);
  assign c1087_inl55 = (((((((((!c962_inl55 && !c964_inl55) && !c966_inl55) && !c968_inl55) && !c970_inl55) && !c972_inl55) && !c974_inl55) && !c976_inl55) && !c978_inl55) && c980_inl55);
  assign c1088_inl55 = ((((((((((!c962_inl55 && !c964_inl55) && !c966_inl55) && !c968_inl55) && !c970_inl55) && !c972_inl55) && !c974_inl55) && !c976_inl55) && !c978_inl55) && !c980_inl55) && c982_inl55);
  assign c1089_inl55 = (((((((((((!c962_inl55 && !c964_inl55) && !c966_inl55) && !c968_inl55) && !c970_inl55) && !c972_inl55) && !c974_inl55) && !c976_inl55) && !c978_inl55) && !c980_inl55) && !c982_inl55) && c984_inl55);
  assign c1090_inl55 = ((((((((((((!c962_inl55 && !c964_inl55) && !c966_inl55) && !c968_inl55) && !c970_inl55) && !c972_inl55) && !c974_inl55) && !c976_inl55) && !c978_inl55) && !c980_inl55) && !c982_inl55) && !c984_inl55) && c986_inl55);
  assign c1091_inl55 = (((((((((((((!c962_inl55 && !c964_inl55) && !c966_inl55) && !c968_inl55) && !c970_inl55) && !c972_inl55) && !c974_inl55) && !c976_inl55) && !c978_inl55) && !c980_inl55) && !c982_inl55) && !c984_inl55) && !c986_inl55) && c988_inl55);
  assign c1092_inl55 = ((((((((((((((!c962_inl55 && !c964_inl55) && !c966_inl55) && !c968_inl55) && !c970_inl55) && !c972_inl55) && !c974_inl55) && !c976_inl55) && !c978_inl55) && !c980_inl55) && !c982_inl55) && !c984_inl55) && !c986_inl55) && !c988_inl55) && c990_inl55);
  assign c1093_inl55 = ((((((((((((((!c962_inl55 && !c964_inl55) && !c966_inl55) && !c968_inl55) && !c970_inl55) && !c972_inl55) && !c974_inl55) && !c976_inl55) && !c978_inl55) && !c980_inl55) && !c982_inl55) && !c984_inl55) && !c986_inl55) && !c988_inl55) && !c990_inl55);
  assign c1094_inl52 = (!c998_inl52 && c1001_inl52);
  assign c1095_inl52 = ((!c998_inl52 && !c1001_inl52) && c1004_inl52);
  assign c1096_inl52 = ((!c998_inl52 && !c1001_inl52) && !c1004_inl52);
  assign c1970 = (c886 && c887);
  assign c1971 = (c886 && c888);
  assign c1972 = (c886 && !c888);
  assign c1973 = (c1971 && c1041);
  assign c1974 = (c1971 && c1042);
  assign c1975 = (c1971 && c1043);
  assign c1976 = (c1971 && c1044);
  assign c1977 = (c1971 && c1045);
  assign c1978 = (c1971 && c1046);
  assign c1979 = (c1971 && c1047);
  assign c1980 = (c1971 && c1048);
  assign c1981 = (c1971 && c1049);
  assign c1982 = (c1971 && c1050);
  assign c1983 = (c1971 && c1051);
  assign c1984 = (c1971 && c1052);
  assign c1985 = (c1971 && c1053);
  assign c1986 = (c1971 && c1054);
  assign c1987 = (c1971 && c1055);
  assign c1988 = (c1971 && c1056);
  assign c1989 = (c1971 && c1057);
  assign c1990 = (c1971 && c1058);
  assign c1991 = (c1971 && c1059);
  assign c1992 = (c1971 && c1060);
  assign c1993 = (c1971 && c1061);
  assign c1994 = (c1971 && c1062);
  assign c1995 = (c1971 && c1063);
  assign c1996 = (c1971 && c1064);
  assign c1997 = (c1971 && c1065);
  assign c1998 = (c1971 && c1066);
  assign c1999 = (c1971 && c1067);
  assign c2000 = (c1971 && c1068);
  assign c2001 = (c1971 && c1069);
  assign c2002 = (c1971 && c1070);
  assign c2004 = (c1973 && c879_inl13);
  assign c2005 = (c1973 && c1036_inl13);
  assign c2006 = (c1973 && c1037_inl13);
  assign c2012 = (c1979 && c872_inl33);
  assign c2013 = (c1979 && c1033_inl33);
  assign c2014 = (c1979 && c1034_inl33);
  assign c2015 = (c1979 && c1035_inl33);
  assign c2016 = (c1980 && c882_inl34);
  assign c2017 = (c1980 && c1038_inl34);
  assign c2018 = (c1980 && c1039_inl34);
  assign c2019 = (c1980 && c1040_inl34);
  assign c2021 = (c1982 && c867_inl35);
  assign c2022 = (c1982 && c1030_inl35);
  assign c2023 = (c1982 && c1031_inl35);
  assign c2024 = (c1982 && c1032_inl35);
  assign c2025 = (c1983 && c862_inl36);
  assign c2026 = (c1983 && c1027_inl36);
  assign c2027 = (c1983 && c1028_inl36);
  assign c2028 = (c1983 && c1029_inl36);
  assign c2029 = (c1984 && c857_inl37);
  assign c2030 = (c1984 && c1024_inl37);
  assign c2031 = (c1984 && c1025_inl37);
  assign c2032 = (c1984 && c1026_inl37);
  assign c2033 = (c1985 && c852_inl38);
  assign c2034 = (c1985 && c1021_inl38);
  assign c2035 = (c1985 && c1022_inl38);
  assign c2036 = (c1985 && c1023_inl38);
  assign c2037 = (c1986 && c848_inl39);
  assign c2038 = (c1986 && c1018_inl39);
  assign c2039 = (c1986 && c1019_inl39);
  assign c2040 = (c1986 && c1020_inl39);
  assign c2041 = (c1987 && c843_inl40);
  assign c2042 = (c1987 && !c843_inl40);
  assign c2046 = (c1991 && c998_inl52);
  assign c2047 = (c1991 && c1094_inl52);
  assign c2048 = (c1991 && c1095_inl52);
  assign c2054 = (c1997 && c845_inl54);
  assign c2055 = (c1997 && !c845_inl54);
  assign c2060 = (c2002 && c927);
  assign c2090 = (c2054 && c846_inl54);
  assign c2091 = (c2054 && !c846_inl54);
  assign c2093 = (c2060 && c930_inl55);
  assign c2120 = (c2093 && c933_inl55);
  assign c2124 = (c2012 && c877_inl33);
  assign c2125 = (c2012 && !c877_inl33);
  assign c2126 = (c2022 && c870_inl35);
  assign c2127 = (c2022 && !c870_inl35);
  assign c2128 = (c2026 && c865_inl36);
  assign c2129 = (c2026 && !c865_inl36);
  assign c2130 = (c2030 && c860_inl37);
  assign c2131 = (c2030 && !c860_inl37);
  assign c2132 = (c2034 && c855_inl38);
  assign c2133 = (c2034 && !c855_inl38);
  assign c2139 = (c2060 && !c930_inl55);
  assign c2140 = (c2093 && !c933_inl55);
  assign c2146 = ((c2041 || c2042) && c924);
  assign c2148 = (((c2139 || c2140) || c2120) && c935_inl55);
  assign c2151 = (c2148 && c938_inl55);
  assign c2152 = (c2148 && !c938_inl55);
  assign c2155 = (c2151 && c939_inl55);
  assign c2156 = (c2151 && !c939_inl55);
  assign c2166 = (((c2139 || c2140) || c2120) && !c935_inl55);
  assign c2167 = ((c2152 || c2155) || c2156);
  assign c2168 = ((c2166 || c2167) && c942_inl55);
  assign c2169 = ((c2166 || c2167) && !c942_inl55);
  assign c2170 = ((c2169 || c2168) && c944_inl55);
  assign c2171 = ((c2169 || c2168) && !c944_inl55);
  assign c2172 = ((c2171 || c2170) && c946_inl55);
  assign c2173 = ((c2171 || c2170) && c1072_inl55);
  assign c2174 = ((c2171 || c2170) && c1073_inl55);
  assign c2175 = ((c2171 || c2170) && c1074_inl55);
  assign c2176 = ((c2171 || c2170) && c1075_inl55);
  assign c2177 = ((c2171 || c2170) && c1076_inl55);
  assign c2178 = ((c2171 || c2170) && c1077_inl55);
  assign c2179 = ((c2171 || c2170) && c1078_inl55);
  assign c2180 = ((((((((c2179 || c2177) || c2176) || c2175) || c2174) || c2173) || c2172) || c2178) && c960_inl55);
  assign c2181 = ((((((((c2179 || c2177) || c2176) || c2175) || c2174) || c2173) || c2172) || c2178) && !c960_inl55);
  assign c2182 = ((c2181 || c2180) && c962_inl55);
  assign c2183 = ((c2181 || c2180) && c1079_inl55);
  assign c2184 = ((c2181 || c2180) && c1080_inl55);
  assign c2185 = ((c2181 || c2180) && c1081_inl55);
  assign c2186 = ((c2181 || c2180) && c1082_inl55);
  assign c2187 = ((c2181 || c2180) && c1083_inl55);
  assign c2188 = ((c2181 || c2180) && c1084_inl55);
  assign c2189 = ((c2181 || c2180) && c1085_inl55);
  assign c2190 = ((c2181 || c2180) && c1086_inl55);
  assign c2191 = ((c2181 || c2180) && c1087_inl55);
  assign c2192 = ((c2181 || c2180) && c1088_inl55);
  assign c2193 = ((c2181 || c2180) && c1089_inl55);
  assign c2194 = ((c2181 || c2180) && c1090_inl55);
  assign c2195 = ((c2181 || c2180) && c1091_inl55);
  assign c2196 = ((c2181 || c2180) && c1092_inl55);
  assign c2197 = ((c2181 || c2180) && c1093_inl55);
  assign c2198 = ((((((((((((((((c2197 || c2185) || c2195) || c2189) || c2194) || c2193) || c2191) || c2192) || c2184) || c2187) || c2190) || c2183) || c2182) || c2196) || c2186) || c2188) && c992_inl55);
  assign c2199 = ((((((((((((((((c2197 || c2185) || c2195) || c2189) || c2194) || c2193) || c2191) || c2192) || c2184) || c2187) || c2190) || c2183) || c2182) || c2196) || c2186) || c2188) && !c992_inl55);
  assign c2200 = (c886 && c920);
  assign c2201 = (c886 && c921);
  assign c3337 = (c886 && c888);
  assign c3338 = (c886 && !c888);
  assign c3339 = (c3337 && c1041);
  assign c3340 = (c3337 && c1042);
  assign c3341 = (c3337 && c1043);
  assign c3342 = (c3337 && c1044);
  assign c3343 = (c3337 && c1045);
  assign c3344 = (c3337 && c1046);
  assign c3345 = (c3337 && c1047);
  assign c3346 = (c3337 && c1048);
  assign c3347 = (c3337 && c1049);
  assign c3348 = (c3337 && c1050);
  assign c3349 = (c3337 && c1051);
  assign c3350 = (c3337 && c1052);
  assign c3351 = (c3337 && c1053);
  assign c3352 = (c3337 && c1054);
  assign c3353 = (c3337 && c1055);
  assign c3354 = (c3337 && c1056);
  assign c3355 = (c3337 && c1057);
  assign c3356 = (c3337 && c1058);
  assign c3357 = (c3337 && c1059);
  assign c3358 = (c3337 && c1060);
  assign c3359 = (c3337 && c1061);
  assign c3360 = (c3337 && c1062);
  assign c3361 = (c3337 && c1063);
  assign c3362 = (c3337 && c1064);
  assign c3363 = (c3337 && c1065);
  assign c3364 = (c3337 && c1066);
  assign c3365 = (c3337 && c1067);
  assign c3366 = (c3337 && c1068);
  assign c3367 = (c3337 && c1069);
  assign c3368 = (c3337 && c1070);
  assign c3369 = (c3339 && c879_inl13);
  assign c3370 = (c3339 && c1036_inl13);
  assign c3371 = (c3339 && c1037_inl13);
  assign c3372 = (c3345 && c872_inl33);
  assign c3373 = (c3345 && c1033_inl33);
  assign c3374 = (c3345 && c1034_inl33);
  assign c3375 = (c3345 && c1035_inl33);
  assign c3376 = (c3346 && c1040_inl34);
  assign c3377 = (c3348 && c867_inl35);
  assign c3378 = (c3348 && c1030_inl35);
  assign c3379 = (c3348 && c1031_inl35);
  assign c3380 = (c3348 && c1032_inl35);
  assign c3381 = (c3349 && c862_inl36);
  assign c3382 = (c3349 && c1027_inl36);
  assign c3383 = (c3349 && c1028_inl36);
  assign c3384 = (c3349 && c1029_inl36);
  assign c3385 = (c3350 && c857_inl37);
  assign c3386 = (c3350 && c1024_inl37);
  assign c3387 = (c3350 && c1025_inl37);
  assign c3388 = (c3350 && c1026_inl37);
  assign c3389 = (c3351 && c852_inl38);
  assign c3390 = (c3351 && c1021_inl38);
  assign c3391 = (c3351 && c1022_inl38);
  assign c3392 = (c3351 && c1023_inl38);
  assign c3393 = (c3352 && c848_inl39);
  assign c3394 = (c3352 && c1018_inl39);
  assign c3395 = (c3352 && c1019_inl39);
  assign c3396 = (c3352 && c1020_inl39);
  assign c3397 = (c3353 && c843_inl40);
  assign c3398 = (c3353 && !c843_inl40);
  assign c3399 = (c3363 && c845_inl54);
  assign c3400 = (c3363 && !c845_inl54);
  assign c3401 = (c3368 && c927);
  assign c3402 = (c3372 && c877_inl33);
  assign c3403 = (c3372 && !c877_inl33);
  assign c3404 = (((c3346 && c882_inl34) || (c3346 && c1038_inl34)) || (c3346 && c1039_inl34));
  assign c3405 = (c3399 && c846_inl54);
  assign c3406 = (c3399 && !c846_inl54);
  assign c3407 = (c3401 && c930_inl55);
  assign c3408 = (c3407 && c933_inl55);
  assign c3409 = (c3401 && !c930_inl55);
  assign c3410 = (c3407 && !c933_inl55);
  assign c3411 = (((c3409 || c3410) || c3408) && c935_inl55);
  assign c3412 = (c3411 && c938_inl55);
  assign c3413 = (c3411 && !c938_inl55);
  assign c3414 = (c3412 && c939_inl55);
  assign c3415 = (c3412 && !c939_inl55);
  assign c3416 = (((c3409 || c3410) || c3408) && !c935_inl55);
  assign c3417 = ((c3413 || c3414) || c3415);
  assign c3418 = ((c3416 || c3417) && c942_inl55);
  assign c3419 = ((c3416 || c3417) && !c942_inl55);
  assign c3420 = ((c3419 || c3418) && c944_inl55);
  assign c3421 = ((c3419 || c3418) && !c944_inl55);
  assign c3422 = ((c3421 || c3420) && c946_inl55);
  assign c3423 = ((c3421 || c3420) && c1072_inl55);
  assign c3424 = ((c3421 || c3420) && c1073_inl55);
  assign c3425 = ((c3421 || c3420) && c1074_inl55);
  assign c3426 = ((c3421 || c3420) && c1075_inl55);
  assign c3427 = ((c3421 || c3420) && c1076_inl55);
  assign c3428 = ((c3421 || c3420) && c1077_inl55);
  assign c3429 = ((c3421 || c3420) && c1078_inl55);
  assign c3430 = ((((((((c3429 || c3427) || c3426) || c3425) || c3424) || c3423) || c3422) || c3428) && c960_inl55);
  assign c3431 = ((((((((c3429 || c3427) || c3426) || c3425) || c3424) || c3423) || c3422) || c3428) && !c960_inl55);
  assign c3432 = ((c3431 || c3430) && c962_inl55);
  assign c3433 = ((c3431 || c3430) && c1079_inl55);
  assign c3434 = ((c3431 || c3430) && c1080_inl55);
  assign c3435 = ((c3431 || c3430) && c1081_inl55);
  assign c3436 = ((c3431 || c3430) && c1082_inl55);
  assign c3437 = ((c3431 || c3430) && c1083_inl55);
  assign c3438 = ((c3431 || c3430) && c1084_inl55);
  assign c3439 = ((c3431 || c3430) && c1085_inl55);
  assign c3440 = ((c3431 || c3430) && c1086_inl55);
  assign c3441 = ((c3431 || c3430) && c1087_inl55);
  assign c3442 = ((c3431 || c3430) && c1088_inl55);
  assign c3443 = ((c3431 || c3430) && c1089_inl55);
  assign c3444 = ((c3431 || c3430) && c1090_inl55);
  assign c3445 = ((c3431 || c3430) && c1091_inl55);
  assign c3446 = ((c3431 || c3430) && c1092_inl55);
  assign c3447 = ((c3431 || c3430) && c1093_inl55);
  assign c3448 = ((((((((((((((((c3447 || c3435) || c3445) || c3439) || c3444) || c3443) || c3441) || c3442) || c3434) || c3437) || c3440) || c3433) || c3432) || c3446) || c3436) || c3438) && c992_inl55);
  assign c3449 = ((((((((((((((((c3447 || c3435) || c3445) || c3439) || c3444) || c3443) || c3441) || c3442) || c3434) || c3437) || c3440) || c3433) || c3432) || c3446) || c3436) || c3438) && !c992_inl55);
  assign c3450 = (c886 && c920);
  assign c843_inl40 = (write_point0_phase2 == 0);
  assign c845_inl54 = (zero_pop_return0_phase2 == 0);
  assign c846_inl54 = (stack0_top2 == 0);
  assign c848_inl39 = (point0_phase2 == 0);
  assign c849_inl39 = (point0_phase2 == 1);
  assign c850_inl39 = (point0_phase2 == 2);
  assign c852_inl38 = (jump_eq0_phase2 == 0);
  assign c853_inl38 = (jump_eq0_phase2 == 1);
  assign c854_inl38 = (jump_eq0_phase2 == 2);
  assign c855_inl38 = (stack0_top2 == jump_eq0_a2);
  assign c857_inl37 = (jump_ne0_phase2 == 0);
  assign c858_inl37 = (jump_ne0_phase2 == 1);
  assign c859_inl37 = (jump_ne0_phase2 == 2);
  assign c860_inl37 = (stack0_top2 != jump_ne0_a2);
  assign c862_inl36 = (jump_le0_phase2 == 0);
  assign c863_inl36 = (jump_le0_phase2 == 1);
  assign c864_inl36 = (jump_le0_phase2 == 2);
  assign c865_inl36 = (stack0_top2 < jump_le0_a2);
  assign c867_inl35 = (jump_ge0_phase2 == 0);
  assign c868_inl35 = (jump_ge0_phase2 == 1);
  assign c869_inl35 = (jump_ge0_phase2 == 2);
  assign c870_inl35 = (stack0_top2 > jump_ge0_a2);
  assign c872_inl33 = (loop0_phase2 == 0);
  assign c873_inl33 = (loop0_phase2 == 1);
  assign c874_inl33 = (loop0_phase2 == 2);
  assign c875_inl33 = (stack0_top10 != 0);
  assign c876_inl33 = (stack0_top10 > -1);
  assign c877_inl33 = (c875_inl33 && c876_inl33);
  assign c879_inl13 = (lit0_phase2 == 0);
  assign c880_inl13 = (lit0_phase2 == 1);
  assign c882_inl34 = (jump0_phase2 == 0);
  assign c883_inl34 = (jump0_phase2 == 1);
  assign c884_inl34 = (jump0_phase2 == 2);
  assign c886 = (ip2 < 268435455);
  assign c887 = (done_flag2 != 0);
  assign c888 = (opcode4 <= 31);
  assign c889 = (opcode4 == 0);
  assign c890 = (opcode4 == 1);
  assign c891 = (opcode4 == 2);
  assign c892 = (opcode4 == 3);
  assign c893 = (opcode4 == 4);
  assign c894 = (opcode4 == 5);
  assign c895 = (opcode4 == 6);
  assign c896 = (opcode4 == 7);
  assign c897 = (opcode4 == 8);
  assign c898 = (opcode4 == 9);
  assign c899 = (opcode4 == 10);
  assign c900 = (opcode4 == 11);
  assign c901 = (opcode4 == 12);
  assign c902 = (opcode4 == 13);
  assign c903 = (opcode4 == 14);
  assign c904 = (opcode4 == 15);
  assign c905 = (opcode4 == 16);
  assign c906 = (opcode4 == 17);
  assign c907 = (opcode4 == 18);
  assign c908 = (opcode4 == 19);
  assign c909 = (opcode4 == 20);
  assign c910 = (opcode4 == 21);
  assign c911 = (opcode4 == 22);
  assign c912 = (opcode4 == 23);
  assign c913 = (opcode4 == 24);
  assign c914 = (opcode4 == 25);
  assign c915 = (opcode4 == 26);
  assign c916 = (opcode4 == 27);
  assign c917 = (opcode4 == 28);
  assign c918 = (opcode4 == 29);
  assign c919 = (opcode4 == 30);
  assign c920 = (wr_flag4 != 0);
  assign c921 = (done_flag13 != 0);
  assign c924 = (exec_result404 != 0);
  assign c927 = (t926 == 0);
  assign c930_inl55 = (t929_inl55 == 1);
  assign c933_inl55 = (t932_inl55 == 13);
  assign c935_inl55 = (t934_inl55 == 1);
  assign c936_inl55 = (stack0_top2 > 0);
  assign c937_inl55 = (stack0_top2 < 128);
  assign c938_inl55 = (c936_inl55 && c937_inl55);
  assign c939_inl55 = (stack0_top2 == 8);
  assign c942_inl55 = (t941_inl55 == 1);
  assign c944_inl55 = (t943_inl55 == 2);
  assign c946_inl55 = (t945_inl55 == -1);
  assign c948_inl55 = (t947_inl55 == -2);
  assign c950_inl55 = (t949_inl55 == -3);
  assign c952_inl55 = (t951_inl55 == -4);
  assign c954_inl55 = (t953_inl55 == -5);
  assign c956_inl55 = (t955_inl55 == -6);
  assign c958_inl55 = (t957_inl55 == -7);
  assign c960_inl55 = (t959_inl55 == -8);
  assign c962_inl55 = (t961_inl55 == -1);
  assign c964_inl55 = (t963_inl55 == -2);
  assign c966_inl55 = (t965_inl55 == -3);
  assign c968_inl55 = (t967_inl55 == -4);
  assign c970_inl55 = (t969_inl55 == -5);
  assign c972_inl55 = (t971_inl55 == -6);
  assign c974_inl55 = (t973_inl55 == -7);
  assign c976_inl55 = (t975_inl55 == -8);
  assign c978_inl55 = (t977_inl55 == -9);
  assign c980_inl55 = (t979_inl55 == -10);
  assign c982_inl55 = (t981_inl55 == -11);
  assign c984_inl55 = (t983_inl55 == -12);
  assign c986_inl55 = (t985_inl55 == -13);
  assign c988_inl55 = (t987_inl55 == -14);
  assign c990_inl55 = (t989_inl55 == -15);
  assign c992_inl55 = (t991_inl55 == 1);
  assign c996_inl52 = (stack0_second2 < 0);
  assign c997_inl52 = (stack0_top2 < 0);
  assign c998_inl52 = (c996_inl52 && c997_inl52);
  assign c999_inl52 = (stack0_second2 > 0);
  assign done_flag13 = (c1971 && c889) ? done_flag2 : ((c2004 || c2005) || c2006) ? exec_result135 : c1974 ? done_flag2 : c1975 ? done_flag2 : c1976 ? done_flag2 : c1977 ? done_flag2 : c1978 ? done_flag2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? exec_result336 : (((c2019 || c2017) || c2018) || c2016) ? exec_result346 : c1981 ? done_flag2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? exec_result357 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? exec_result367 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? exec_result377 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? exec_result387 : (((c2038 || c2040) || c2037) || c2039) ? exec_result396 : (c2041 || c2042) ? exec_result404 : c1988 ? done_flag2 : c1989 ? done_flag2 : c1990 ? done_flag2 : c1991 ? done_flag2 : c1992 ? done_flag2 : c1993 ? done_flag2 : c1994 ? done_flag2 : c1995 ? done_flag2 : c1996 ? done_flag2 : ((c2055 || c2091) || c2090) ? exec_result545 : c1998 ? done_flag2 : c1999 ? done_flag2 : c2000 ? done_flag2 : c2001 ? done_flag2 : (c2199 || c2198) ? done_flag2 : (c2002 && !c927) ? done_flag2 : c1972 ? done_flag2 : 'bz;
  assign exec_result135 = c2004 ? 0 : c2005 ? 0 : c2006 ? 1 : 'bz;
  assign exec_result346 = c2016 ? 0 : c2017 ? 0 : c2018 ? 0 : c2019 ? 1 : 'bz;
  assign exec_result357 = c2021 ? 0 : c2022 ? t2771 : c2023 ? 0 : c2024 ? 1 : 'bz;
  assign exec_result367 = c2025 ? 0 : c2026 ? t2778 : c2027 ? 0 : c2028 ? 1 : 'bz;
  assign exec_result377 = c2029 ? 0 : c2030 ? t2785 : c2031 ? 0 : c2032 ? 1 : 'bz;
  assign exec_result387 = c2033 ? 0 : c2034 ? t2792 : c2035 ? 0 : c2036 ? 1 : 'bz;
  assign exec_result396 = c2037 ? 0 : c2038 ? 0 : c2039 ? 0 : c2040 ? 1 : 'bz;
  assign exec_result404 = c2041 ? 0 : c2042 ? 1 : 'bz;
  assign exec_result545 = c2090 ? 0 : c2091 ? 1 : c2055 ? 1 : 'bz;
  assign ip15 = (t928 - 1);
  assign ip16 = (c1971 && c889) ? ip2 : ((c2004 || c2005) || c2006) ? lit0_ip4 : c1974 ? ip2 : c1975 ? ip2 : c1976 ? ip2 : c1977 ? ip2 : c1978 ? ip2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? loop0_ip5 : (((c2019 || c2017) || c2018) || c2016) ? jump0_ip5 : c1981 ? address0_top2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? jump_ge0_ip5 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? jump_le0_ip5 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? jump_ne0_ip5 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? jump_eq0_ip5 : (((c2038 || c2040) || c2037) || c2039) ? point0_ip5 : (c2041 || c2042) ? write_point0_ip4 : c1988 ? ip2 : c1989 ? ip2 : c1990 ? ip2 : c1991 ? ip2 : c1992 ? ip2 : c1993 ? ip2 : c1994 ? ip2 : c1995 ? ip2 : c1996 ? ip2 : ((c2055 || c2091) || c2090) ? zero_pop_return0_ip5 : c1998 ? ip2 : c1999 ? ip2 : c2000 ? ip2 : c2001 ? ip2 : (c2199 || c2198) ? ip_inl554 : (c2002 && !c927) ? ip2 : c1972 ? ip15 : 'bz;
  assign ip17 = (ip16 + 1);
  assign ip18 = c2201 ? ip17 : (c886 && !c921) ? ip16 : 'bz;
  assign ip_inl554 = c2182 ? ip2 : c2183 ? ip2 : c2184 ? ip2 : c2185 ? ip2 : c2186 ? ip2 : c2187 ? ip2 : c2188 ? ip2 : c2189 ? ip2 : c2190 ? 268435455 : c2191 ? ip2 : c2192 ? ip2 : c2193 ? ip2 : c2194 ? ip2 : c2195 ? ip2 : c2196 ? ip2 : ((c2181 || c2180) && c1093_inl55) ? ip2 : 'bz;
  assign jump0_ip3 = (ip2 + 1);
  assign jump0_ip4 = (mem_data - 1);
  assign jump0_ip5 = c2016 ? jump0_ip3 : c2017 ? jump0_ip2 : c2018 ? jump0_ip4 : c2019 ? jump0_ip2 : 'bz;
  assign jump0_ip6 = (c1971 && c889) ? jump0_ip2 : ((c2004 || c2005) || c2006) ? jump0_ip2 : c1974 ? jump0_ip2 : c1975 ? jump0_ip2 : c1976 ? jump0_ip2 : c1977 ? jump0_ip2 : c1978 ? jump0_ip2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? jump0_ip2 : (((c2019 || c2017) || c2018) || c2016) ? jump0_ip5 : c1981 ? jump0_ip2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? jump0_ip2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? jump0_ip2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? jump0_ip2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? jump0_ip2 : (((c2038 || c2040) || c2037) || c2039) ? jump0_ip2 : (c2041 || c2042) ? jump0_ip2 : c1988 ? jump0_ip2 : c1989 ? jump0_ip2 : c1990 ? jump0_ip2 : c1991 ? jump0_ip2 : c1992 ? jump0_ip2 : c1993 ? jump0_ip2 : c1994 ? jump0_ip2 : c1995 ? jump0_ip2 : c1996 ? jump0_ip2 : ((c2055 || c2091) || c2090) ? jump0_ip2 : c1998 ? jump0_ip2 : c1999 ? jump0_ip2 : c2000 ? jump0_ip2 : c2001 ? jump0_ip2 : (c2199 || c2198) ? jump0_ip2 : (c2002 && !c927) ? jump0_ip2 : c1972 ? jump0_ip2 : 'bz;
  assign jump0_phase7 = c2016 ? 1 : c2017 ? 2 : c2018 ? 3 : c2019 ? 0 : 'bz;
  assign jump0_phase8 = (c1971 && c889) ? jump0_phase2 : ((c2004 || c2005) || c2006) ? jump0_phase2 : c1974 ? jump0_phase2 : c1975 ? jump0_phase2 : c1976 ? jump0_phase2 : c1977 ? jump0_phase2 : c1978 ? jump0_phase2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? jump0_phase2 : (((c2019 || c2017) || c2018) || c2016) ? jump0_phase7 : c1981 ? jump0_phase2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? jump0_phase2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? jump0_phase2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? jump0_phase2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? jump0_phase2 : (((c2038 || c2040) || c2037) || c2039) ? jump0_phase2 : (c2041 || c2042) ? jump0_phase2 : c1988 ? jump0_phase2 : c1989 ? jump0_phase2 : c1990 ? jump0_phase2 : c1991 ? jump0_phase2 : c1992 ? jump0_phase2 : c1993 ? jump0_phase2 : c1994 ? jump0_phase2 : c1995 ? jump0_phase2 : c1996 ? jump0_phase2 : ((c2055 || c2091) || c2090) ? jump0_phase2 : c1998 ? jump0_phase2 : c1999 ? jump0_phase2 : c2000 ? jump0_phase2 : c2001 ? jump0_phase2 : (c2199 || c2198) ? jump0_phase2 : (c2002 && !c927) ? jump0_phase2 : c1972 ? jump0_phase2 : 'bz;
  assign jump_eq0_a4 = c2033 ? stack0_top2 : c2034 ? jump_eq0_a2 : c2035 ? jump_eq0_a2 : c2036 ? jump_eq0_a2 : 'bz;
  assign jump_eq0_a5 = (c1971 && c889) ? jump_eq0_a2 : ((c2004 || c2005) || c2006) ? jump_eq0_a2 : c1974 ? jump_eq0_a2 : c1975 ? jump_eq0_a2 : c1976 ? jump_eq0_a2 : c1977 ? jump_eq0_a2 : c1978 ? jump_eq0_a2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? jump_eq0_a2 : (((c2019 || c2017) || c2018) || c2016) ? jump_eq0_a2 : c1981 ? jump_eq0_a2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? jump_eq0_a2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? jump_eq0_a2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? jump_eq0_a2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? jump_eq0_a4 : (((c2038 || c2040) || c2037) || c2039) ? jump_eq0_a2 : (c2041 || c2042) ? jump_eq0_a2 : c1988 ? jump_eq0_a2 : c1989 ? jump_eq0_a2 : c1990 ? jump_eq0_a2 : c1991 ? jump_eq0_a2 : c1992 ? jump_eq0_a2 : c1993 ? jump_eq0_a2 : c1994 ? jump_eq0_a2 : c1995 ? jump_eq0_a2 : c1996 ? jump_eq0_a2 : ((c2055 || c2091) || c2090) ? jump_eq0_a2 : c1998 ? jump_eq0_a2 : c1999 ? jump_eq0_a2 : c2000 ? jump_eq0_a2 : c2001 ? jump_eq0_a2 : (c2199 || c2198) ? jump_eq0_a2 : (c2002 && !c927) ? jump_eq0_a2 : c1972 ? jump_eq0_a2 : 'bz;
  assign jump_eq0_ip3 = (ip2 + 1);
  assign jump_eq0_ip4 = (mem_data - 1);
  assign jump_eq0_ip5 = c2033 ? jump_eq0_ip3 : c2034 ? jump_eq0_ip2 : c2035 ? jump_eq0_ip4 : c2036 ? jump_eq0_ip2 : 'bz;
  assign jump_eq0_ip6 = (c1971 && c889) ? jump_eq0_ip2 : ((c2004 || c2005) || c2006) ? jump_eq0_ip2 : c1974 ? jump_eq0_ip2 : c1975 ? jump_eq0_ip2 : c1976 ? jump_eq0_ip2 : c1977 ? jump_eq0_ip2 : c1978 ? jump_eq0_ip2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? jump_eq0_ip2 : (((c2019 || c2017) || c2018) || c2016) ? jump_eq0_ip2 : c1981 ? jump_eq0_ip2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? jump_eq0_ip2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? jump_eq0_ip2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? jump_eq0_ip2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? jump_eq0_ip5 : (((c2038 || c2040) || c2037) || c2039) ? jump_eq0_ip2 : (c2041 || c2042) ? jump_eq0_ip2 : c1988 ? jump_eq0_ip2 : c1989 ? jump_eq0_ip2 : c1990 ? jump_eq0_ip2 : c1991 ? jump_eq0_ip2 : c1992 ? jump_eq0_ip2 : c1993 ? jump_eq0_ip2 : c1994 ? jump_eq0_ip2 : c1995 ? jump_eq0_ip2 : c1996 ? jump_eq0_ip2 : ((c2055 || c2091) || c2090) ? jump_eq0_ip2 : c1998 ? jump_eq0_ip2 : c1999 ? jump_eq0_ip2 : c2000 ? jump_eq0_ip2 : c2001 ? jump_eq0_ip2 : (c2199 || c2198) ? jump_eq0_ip2 : (c2002 && !c927) ? jump_eq0_ip2 : c1972 ? jump_eq0_ip2 : 'bz;
  assign jump_eq0_phase8 = c2033 ? 1 : c2034 ? t2795 : c2035 ? 3 : c2036 ? 0 : 'bz;
  assign jump_eq0_phase9 = (c1971 && c889) ? jump_eq0_phase2 : ((c2004 || c2005) || c2006) ? jump_eq0_phase2 : c1974 ? jump_eq0_phase2 : c1975 ? jump_eq0_phase2 : c1976 ? jump_eq0_phase2 : c1977 ? jump_eq0_phase2 : c1978 ? jump_eq0_phase2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? jump_eq0_phase2 : (((c2019 || c2017) || c2018) || c2016) ? jump_eq0_phase2 : c1981 ? jump_eq0_phase2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? jump_eq0_phase2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? jump_eq0_phase2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? jump_eq0_phase2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? jump_eq0_phase8 : (((c2038 || c2040) || c2037) || c2039) ? jump_eq0_phase2 : (c2041 || c2042) ? jump_eq0_phase2 : c1988 ? jump_eq0_phase2 : c1989 ? jump_eq0_phase2 : c1990 ? jump_eq0_phase2 : c1991 ? jump_eq0_phase2 : c1992 ? jump_eq0_phase2 : c1993 ? jump_eq0_phase2 : c1994 ? jump_eq0_phase2 : c1995 ? jump_eq0_phase2 : c1996 ? jump_eq0_phase2 : ((c2055 || c2091) || c2090) ? jump_eq0_phase2 : c1998 ? jump_eq0_phase2 : c1999 ? jump_eq0_phase2 : c2000 ? jump_eq0_phase2 : c2001 ? jump_eq0_phase2 : (c2199 || c2198) ? jump_eq0_phase2 : (c2002 && !c927) ? jump_eq0_phase2 : c1972 ? jump_eq0_phase2 : 'bz;
  assign jump_ge0_a4 = c2021 ? stack0_top2 : c2022 ? jump_ge0_a2 : c2023 ? jump_ge0_a2 : c2024 ? jump_ge0_a2 : 'bz;
  assign jump_ge0_a5 = (c1971 && c889) ? jump_ge0_a2 : ((c2004 || c2005) || c2006) ? jump_ge0_a2 : c1974 ? jump_ge0_a2 : c1975 ? jump_ge0_a2 : c1976 ? jump_ge0_a2 : c1977 ? jump_ge0_a2 : c1978 ? jump_ge0_a2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? jump_ge0_a2 : (((c2019 || c2017) || c2018) || c2016) ? jump_ge0_a2 : c1981 ? jump_ge0_a2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? jump_ge0_a4 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? jump_ge0_a2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? jump_ge0_a2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? jump_ge0_a2 : (((c2038 || c2040) || c2037) || c2039) ? jump_ge0_a2 : (c2041 || c2042) ? jump_ge0_a2 : c1988 ? jump_ge0_a2 : c1989 ? jump_ge0_a2 : c1990 ? jump_ge0_a2 : c1991 ? jump_ge0_a2 : c1992 ? jump_ge0_a2 : c1993 ? jump_ge0_a2 : c1994 ? jump_ge0_a2 : c1995 ? jump_ge0_a2 : c1996 ? jump_ge0_a2 : ((c2055 || c2091) || c2090) ? jump_ge0_a2 : c1998 ? jump_ge0_a2 : c1999 ? jump_ge0_a2 : c2000 ? jump_ge0_a2 : c2001 ? jump_ge0_a2 : (c2199 || c2198) ? jump_ge0_a2 : (c2002 && !c927) ? jump_ge0_a2 : c1972 ? jump_ge0_a2 : 'bz;
  assign jump_ge0_ip3 = (ip2 + 1);
  assign jump_ge0_ip4 = (mem_data - 1);
  assign jump_ge0_ip5 = c2021 ? jump_ge0_ip3 : c2022 ? jump_ge0_ip2 : c2023 ? jump_ge0_ip4 : c2024 ? jump_ge0_ip2 : 'bz;
  assign jump_ge0_ip6 = (c1971 && c889) ? jump_ge0_ip2 : ((c2004 || c2005) || c2006) ? jump_ge0_ip2 : c1974 ? jump_ge0_ip2 : c1975 ? jump_ge0_ip2 : c1976 ? jump_ge0_ip2 : c1977 ? jump_ge0_ip2 : c1978 ? jump_ge0_ip2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? jump_ge0_ip2 : (((c2019 || c2017) || c2018) || c2016) ? jump_ge0_ip2 : c1981 ? jump_ge0_ip2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? jump_ge0_ip5 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? jump_ge0_ip2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? jump_ge0_ip2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? jump_ge0_ip2 : (((c2038 || c2040) || c2037) || c2039) ? jump_ge0_ip2 : (c2041 || c2042) ? jump_ge0_ip2 : c1988 ? jump_ge0_ip2 : c1989 ? jump_ge0_ip2 : c1990 ? jump_ge0_ip2 : c1991 ? jump_ge0_ip2 : c1992 ? jump_ge0_ip2 : c1993 ? jump_ge0_ip2 : c1994 ? jump_ge0_ip2 : c1995 ? jump_ge0_ip2 : c1996 ? jump_ge0_ip2 : ((c2055 || c2091) || c2090) ? jump_ge0_ip2 : c1998 ? jump_ge0_ip2 : c1999 ? jump_ge0_ip2 : c2000 ? jump_ge0_ip2 : c2001 ? jump_ge0_ip2 : (c2199 || c2198) ? jump_ge0_ip2 : (c2002 && !c927) ? jump_ge0_ip2 : c1972 ? jump_ge0_ip2 : 'bz;
  assign jump_ge0_phase8 = c2021 ? 1 : c2022 ? t2774 : c2023 ? 3 : c2024 ? 0 : 'bz;
  assign jump_ge0_phase9 = (c1971 && c889) ? jump_ge0_phase2 : ((c2004 || c2005) || c2006) ? jump_ge0_phase2 : c1974 ? jump_ge0_phase2 : c1975 ? jump_ge0_phase2 : c1976 ? jump_ge0_phase2 : c1977 ? jump_ge0_phase2 : c1978 ? jump_ge0_phase2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? jump_ge0_phase2 : (((c2019 || c2017) || c2018) || c2016) ? jump_ge0_phase2 : c1981 ? jump_ge0_phase2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? jump_ge0_phase8 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? jump_ge0_phase2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? jump_ge0_phase2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? jump_ge0_phase2 : (((c2038 || c2040) || c2037) || c2039) ? jump_ge0_phase2 : (c2041 || c2042) ? jump_ge0_phase2 : c1988 ? jump_ge0_phase2 : c1989 ? jump_ge0_phase2 : c1990 ? jump_ge0_phase2 : c1991 ? jump_ge0_phase2 : c1992 ? jump_ge0_phase2 : c1993 ? jump_ge0_phase2 : c1994 ? jump_ge0_phase2 : c1995 ? jump_ge0_phase2 : c1996 ? jump_ge0_phase2 : ((c2055 || c2091) || c2090) ? jump_ge0_phase2 : c1998 ? jump_ge0_phase2 : c1999 ? jump_ge0_phase2 : c2000 ? jump_ge0_phase2 : c2001 ? jump_ge0_phase2 : (c2199 || c2198) ? jump_ge0_phase2 : (c2002 && !c927) ? jump_ge0_phase2 : c1972 ? jump_ge0_phase2 : 'bz;
  assign jump_le0_a4 = c2025 ? stack0_top2 : c2026 ? jump_le0_a2 : c2027 ? jump_le0_a2 : c2028 ? jump_le0_a2 : 'bz;
  assign jump_le0_a5 = (c1971 && c889) ? jump_le0_a2 : ((c2004 || c2005) || c2006) ? jump_le0_a2 : c1974 ? jump_le0_a2 : c1975 ? jump_le0_a2 : c1976 ? jump_le0_a2 : c1977 ? jump_le0_a2 : c1978 ? jump_le0_a2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? jump_le0_a2 : (((c2019 || c2017) || c2018) || c2016) ? jump_le0_a2 : c1981 ? jump_le0_a2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? jump_le0_a2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? jump_le0_a4 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? jump_le0_a2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? jump_le0_a2 : (((c2038 || c2040) || c2037) || c2039) ? jump_le0_a2 : (c2041 || c2042) ? jump_le0_a2 : c1988 ? jump_le0_a2 : c1989 ? jump_le0_a2 : c1990 ? jump_le0_a2 : c1991 ? jump_le0_a2 : c1992 ? jump_le0_a2 : c1993 ? jump_le0_a2 : c1994 ? jump_le0_a2 : c1995 ? jump_le0_a2 : c1996 ? jump_le0_a2 : ((c2055 || c2091) || c2090) ? jump_le0_a2 : c1998 ? jump_le0_a2 : c1999 ? jump_le0_a2 : c2000 ? jump_le0_a2 : c2001 ? jump_le0_a2 : (c2199 || c2198) ? jump_le0_a2 : (c2002 && !c927) ? jump_le0_a2 : c1972 ? jump_le0_a2 : 'bz;
  assign jump_le0_ip3 = (ip2 + 1);
  assign jump_le0_ip4 = (mem_data - 1);
  assign jump_le0_ip5 = c2025 ? jump_le0_ip3 : c2026 ? jump_le0_ip2 : c2027 ? jump_le0_ip4 : c2028 ? jump_le0_ip2 : 'bz;
  assign jump_le0_ip6 = (c1971 && c889) ? jump_le0_ip2 : ((c2004 || c2005) || c2006) ? jump_le0_ip2 : c1974 ? jump_le0_ip2 : c1975 ? jump_le0_ip2 : c1976 ? jump_le0_ip2 : c1977 ? jump_le0_ip2 : c1978 ? jump_le0_ip2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? jump_le0_ip2 : (((c2019 || c2017) || c2018) || c2016) ? jump_le0_ip2 : c1981 ? jump_le0_ip2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? jump_le0_ip2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? jump_le0_ip5 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? jump_le0_ip2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? jump_le0_ip2 : (((c2038 || c2040) || c2037) || c2039) ? jump_le0_ip2 : (c2041 || c2042) ? jump_le0_ip2 : c1988 ? jump_le0_ip2 : c1989 ? jump_le0_ip2 : c1990 ? jump_le0_ip2 : c1991 ? jump_le0_ip2 : c1992 ? jump_le0_ip2 : c1993 ? jump_le0_ip2 : c1994 ? jump_le0_ip2 : c1995 ? jump_le0_ip2 : c1996 ? jump_le0_ip2 : ((c2055 || c2091) || c2090) ? jump_le0_ip2 : c1998 ? jump_le0_ip2 : c1999 ? jump_le0_ip2 : c2000 ? jump_le0_ip2 : c2001 ? jump_le0_ip2 : (c2199 || c2198) ? jump_le0_ip2 : (c2002 && !c927) ? jump_le0_ip2 : c1972 ? jump_le0_ip2 : 'bz;
  assign jump_le0_phase8 = c2025 ? 1 : c2026 ? t2781 : c2027 ? 3 : c2028 ? 0 : 'bz;
  assign jump_le0_phase9 = (c1971 && c889) ? jump_le0_phase2 : ((c2004 || c2005) || c2006) ? jump_le0_phase2 : c1974 ? jump_le0_phase2 : c1975 ? jump_le0_phase2 : c1976 ? jump_le0_phase2 : c1977 ? jump_le0_phase2 : c1978 ? jump_le0_phase2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? jump_le0_phase2 : (((c2019 || c2017) || c2018) || c2016) ? jump_le0_phase2 : c1981 ? jump_le0_phase2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? jump_le0_phase2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? jump_le0_phase8 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? jump_le0_phase2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? jump_le0_phase2 : (((c2038 || c2040) || c2037) || c2039) ? jump_le0_phase2 : (c2041 || c2042) ? jump_le0_phase2 : c1988 ? jump_le0_phase2 : c1989 ? jump_le0_phase2 : c1990 ? jump_le0_phase2 : c1991 ? jump_le0_phase2 : c1992 ? jump_le0_phase2 : c1993 ? jump_le0_phase2 : c1994 ? jump_le0_phase2 : c1995 ? jump_le0_phase2 : c1996 ? jump_le0_phase2 : ((c2055 || c2091) || c2090) ? jump_le0_phase2 : c1998 ? jump_le0_phase2 : c1999 ? jump_le0_phase2 : c2000 ? jump_le0_phase2 : c2001 ? jump_le0_phase2 : (c2199 || c2198) ? jump_le0_phase2 : (c2002 && !c927) ? jump_le0_phase2 : c1972 ? jump_le0_phase2 : 'bz;
  assign jump_ne0_a4 = c2029 ? stack0_top2 : c2030 ? jump_ne0_a2 : c2031 ? jump_ne0_a2 : c2032 ? jump_ne0_a2 : 'bz;
  assign jump_ne0_a5 = (c1971 && c889) ? jump_ne0_a2 : ((c2004 || c2005) || c2006) ? jump_ne0_a2 : c1974 ? jump_ne0_a2 : c1975 ? jump_ne0_a2 : c1976 ? jump_ne0_a2 : c1977 ? jump_ne0_a2 : c1978 ? jump_ne0_a2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? jump_ne0_a2 : (((c2019 || c2017) || c2018) || c2016) ? jump_ne0_a2 : c1981 ? jump_ne0_a2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? jump_ne0_a2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? jump_ne0_a2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? jump_ne0_a4 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? jump_ne0_a2 : (((c2038 || c2040) || c2037) || c2039) ? jump_ne0_a2 : (c2041 || c2042) ? jump_ne0_a2 : c1988 ? jump_ne0_a2 : c1989 ? jump_ne0_a2 : c1990 ? jump_ne0_a2 : c1991 ? jump_ne0_a2 : c1992 ? jump_ne0_a2 : c1993 ? jump_ne0_a2 : c1994 ? jump_ne0_a2 : c1995 ? jump_ne0_a2 : c1996 ? jump_ne0_a2 : ((c2055 || c2091) || c2090) ? jump_ne0_a2 : c1998 ? jump_ne0_a2 : c1999 ? jump_ne0_a2 : c2000 ? jump_ne0_a2 : c2001 ? jump_ne0_a2 : (c2199 || c2198) ? jump_ne0_a2 : (c2002 && !c927) ? jump_ne0_a2 : c1972 ? jump_ne0_a2 : 'bz;
  assign jump_ne0_ip3 = (ip2 + 1);
  assign jump_ne0_ip4 = (mem_data - 1);
  assign jump_ne0_ip5 = c2029 ? jump_ne0_ip3 : c2030 ? jump_ne0_ip2 : c2031 ? jump_ne0_ip4 : c2032 ? jump_ne0_ip2 : 'bz;
  assign jump_ne0_ip6 = (c1971 && c889) ? jump_ne0_ip2 : ((c2004 || c2005) || c2006) ? jump_ne0_ip2 : c1974 ? jump_ne0_ip2 : c1975 ? jump_ne0_ip2 : c1976 ? jump_ne0_ip2 : c1977 ? jump_ne0_ip2 : c1978 ? jump_ne0_ip2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? jump_ne0_ip2 : (((c2019 || c2017) || c2018) || c2016) ? jump_ne0_ip2 : c1981 ? jump_ne0_ip2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? jump_ne0_ip2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? jump_ne0_ip2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? jump_ne0_ip5 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? jump_ne0_ip2 : (((c2038 || c2040) || c2037) || c2039) ? jump_ne0_ip2 : (c2041 || c2042) ? jump_ne0_ip2 : c1988 ? jump_ne0_ip2 : c1989 ? jump_ne0_ip2 : c1990 ? jump_ne0_ip2 : c1991 ? jump_ne0_ip2 : c1992 ? jump_ne0_ip2 : c1993 ? jump_ne0_ip2 : c1994 ? jump_ne0_ip2 : c1995 ? jump_ne0_ip2 : c1996 ? jump_ne0_ip2 : ((c2055 || c2091) || c2090) ? jump_ne0_ip2 : c1998 ? jump_ne0_ip2 : c1999 ? jump_ne0_ip2 : c2000 ? jump_ne0_ip2 : c2001 ? jump_ne0_ip2 : (c2199 || c2198) ? jump_ne0_ip2 : (c2002 && !c927) ? jump_ne0_ip2 : c1972 ? jump_ne0_ip2 : 'bz;
  assign jump_ne0_phase8 = c2029 ? 1 : c2030 ? t2788 : c2031 ? 3 : c2032 ? 0 : 'bz;
  assign jump_ne0_phase9 = (c1971 && c889) ? jump_ne0_phase2 : ((c2004 || c2005) || c2006) ? jump_ne0_phase2 : c1974 ? jump_ne0_phase2 : c1975 ? jump_ne0_phase2 : c1976 ? jump_ne0_phase2 : c1977 ? jump_ne0_phase2 : c1978 ? jump_ne0_phase2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? jump_ne0_phase2 : (((c2019 || c2017) || c2018) || c2016) ? jump_ne0_phase2 : c1981 ? jump_ne0_phase2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? jump_ne0_phase2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? jump_ne0_phase2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? jump_ne0_phase8 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? jump_ne0_phase2 : (((c2038 || c2040) || c2037) || c2039) ? jump_ne0_phase2 : (c2041 || c2042) ? jump_ne0_phase2 : c1988 ? jump_ne0_phase2 : c1989 ? jump_ne0_phase2 : c1990 ? jump_ne0_phase2 : c1991 ? jump_ne0_phase2 : c1992 ? jump_ne0_phase2 : c1993 ? jump_ne0_phase2 : c1994 ? jump_ne0_phase2 : c1995 ? jump_ne0_phase2 : c1996 ? jump_ne0_phase2 : ((c2055 || c2091) || c2090) ? jump_ne0_phase2 : c1998 ? jump_ne0_phase2 : c1999 ? jump_ne0_phase2 : c2000 ? jump_ne0_phase2 : c2001 ? jump_ne0_phase2 : (c2199 || c2198) ? jump_ne0_phase2 : (c2002 && !c927) ? jump_ne0_phase2 : c1972 ? jump_ne0_phase2 : 'bz;
  assign lit0_ip3 = (ip2 + 1);
  assign lit0_ip4 = c2004 ? lit0_ip3 : c2005 ? lit0_ip2 : c2006 ? lit0_ip2 : 'bz;
  assign lit0_ip5 = (c1971 && c889) ? lit0_ip2 : ((c2004 || c2005) || c2006) ? lit0_ip4 : c1974 ? lit0_ip2 : c1975 ? lit0_ip2 : c1976 ? lit0_ip2 : c1977 ? lit0_ip2 : c1978 ? lit0_ip2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? lit0_ip2 : (((c2019 || c2017) || c2018) || c2016) ? lit0_ip2 : c1981 ? lit0_ip2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? lit0_ip2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? lit0_ip2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? lit0_ip2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? lit0_ip2 : (((c2038 || c2040) || c2037) || c2039) ? lit0_ip2 : (c2041 || c2042) ? lit0_ip2 : c1988 ? lit0_ip2 : c1989 ? lit0_ip2 : c1990 ? lit0_ip2 : c1991 ? lit0_ip2 : c1992 ? lit0_ip2 : c1993 ? lit0_ip2 : c1994 ? lit0_ip2 : c1995 ? lit0_ip2 : c1996 ? lit0_ip2 : ((c2055 || c2091) || c2090) ? lit0_ip2 : c1998 ? lit0_ip2 : c1999 ? lit0_ip2 : c2000 ? lit0_ip2 : c2001 ? lit0_ip2 : (c2199 || c2198) ? lit0_ip2 : (c2002 && !c927) ? lit0_ip2 : c1972 ? lit0_ip2 : 'bz;
  assign lit0_phase6 = c2004 ? 1 : c2005 ? 2 : c2006 ? 0 : 'bz;
  assign lit0_phase7 = (c1971 && c889) ? lit0_phase2 : ((c2004 || c2005) || c2006) ? lit0_phase6 : c1974 ? lit0_phase2 : c1975 ? lit0_phase2 : c1976 ? lit0_phase2 : c1977 ? lit0_phase2 : c1978 ? lit0_phase2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? lit0_phase2 : (((c2019 || c2017) || c2018) || c2016) ? lit0_phase2 : c1981 ? lit0_phase2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? lit0_phase2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? lit0_phase2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? lit0_phase2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? lit0_phase2 : (((c2038 || c2040) || c2037) || c2039) ? lit0_phase2 : (c2041 || c2042) ? lit0_phase2 : c1988 ? lit0_phase2 : c1989 ? lit0_phase2 : c1990 ? lit0_phase2 : c1991 ? lit0_phase2 : c1992 ? lit0_phase2 : c1993 ? lit0_phase2 : c1994 ? lit0_phase2 : c1995 ? lit0_phase2 : c1996 ? lit0_phase2 : ((c2055 || c2091) || c2090) ? lit0_phase2 : c1998 ? lit0_phase2 : c1999 ? lit0_phase2 : c2000 ? lit0_phase2 : c2001 ? lit0_phase2 : (c2199 || c2198) ? lit0_phase2 : (c2002 && !c927) ? lit0_phase2 : c1972 ? lit0_phase2 : 'bz;
  assign loop0_ip3 = (ip2 + 1);
  assign loop0_ip4 = (mem_data - 1);
  assign loop0_ip5 = c2124 ? loop0_ip3 : c2125 ? loop0_ip3 : c2013 ? loop0_ip2 : c2014 ? loop0_ip4 : c2015 ? loop0_ip2 : 'bz;
  assign loop0_ip6 = (c1971 && c889) ? loop0_ip2 : ((c2004 || c2005) || c2006) ? loop0_ip2 : c1974 ? loop0_ip2 : c1975 ? loop0_ip2 : c1976 ? loop0_ip2 : c1977 ? loop0_ip2 : c1978 ? loop0_ip2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? loop0_ip5 : (((c2019 || c2017) || c2018) || c2016) ? loop0_ip2 : c1981 ? loop0_ip2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? loop0_ip2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? loop0_ip2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? loop0_ip2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? loop0_ip2 : (((c2038 || c2040) || c2037) || c2039) ? loop0_ip2 : (c2041 || c2042) ? loop0_ip2 : c1988 ? loop0_ip2 : c1989 ? loop0_ip2 : c1990 ? loop0_ip2 : c1991 ? loop0_ip2 : c1992 ? loop0_ip2 : c1993 ? loop0_ip2 : c1994 ? loop0_ip2 : c1995 ? loop0_ip2 : c1996 ? loop0_ip2 : ((c2055 || c2091) || c2090) ? loop0_ip2 : c1998 ? loop0_ip2 : c1999 ? loop0_ip2 : c2000 ? loop0_ip2 : c2001 ? loop0_ip2 : (c2199 || c2198) ? loop0_ip2 : (c2002 && !c927) ? loop0_ip2 : c1972 ? loop0_ip2 : 'bz;
  assign loop0_phase8 = c2124 ? 1 : c2125 ? 0 : c2013 ? 2 : c2014 ? 3 : c2015 ? 0 : 'bz;
  assign loop0_phase9 = (c1971 && c889) ? loop0_phase2 : ((c2004 || c2005) || c2006) ? loop0_phase2 : c1974 ? loop0_phase2 : c1975 ? loop0_phase2 : c1976 ? loop0_phase2 : c1977 ? loop0_phase2 : c1978 ? loop0_phase2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? loop0_phase8 : (((c2019 || c2017) || c2018) || c2016) ? loop0_phase2 : c1981 ? loop0_phase2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? loop0_phase2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? loop0_phase2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? loop0_phase2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? loop0_phase2 : (((c2038 || c2040) || c2037) || c2039) ? loop0_phase2 : (c2041 || c2042) ? loop0_phase2 : c1988 ? loop0_phase2 : c1989 ? loop0_phase2 : c1990 ? loop0_phase2 : c1991 ? loop0_phase2 : c1992 ? loop0_phase2 : c1993 ? loop0_phase2 : c1994 ? loop0_phase2 : c1995 ? loop0_phase2 : c1996 ? loop0_phase2 : ((c2055 || c2091) || c2090) ? loop0_phase2 : c1998 ? loop0_phase2 : c1999 ? loop0_phase2 : c2000 ? loop0_phase2 : c2001 ? loop0_phase2 : (c2199 || c2198) ? loop0_phase2 : (c2002 && !c927) ? loop0_phase2 : c1972 ? loop0_phase2 : 'bz;
  assign opcode4 = c1970 ? mem_data : (c886 && !c887) ? opcode2 : 'bz;
  assign point0_ip5 = c2037 ? stack0_top2 : c2038 ? point0_ip2 : c2039 ? point0_ip_saved2 : c2040 ? point0_ip2 : 'bz;
  assign point0_ip6 = (c1971 && c889) ? point0_ip2 : ((c2004 || c2005) || c2006) ? point0_ip2 : c1974 ? point0_ip2 : c1975 ? point0_ip2 : c1976 ? point0_ip2 : c1977 ? point0_ip2 : c1978 ? point0_ip2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? point0_ip2 : (((c2019 || c2017) || c2018) || c2016) ? point0_ip2 : c1981 ? point0_ip2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? point0_ip2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? point0_ip2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? point0_ip2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? point0_ip2 : (((c2038 || c2040) || c2037) || c2039) ? point0_ip5 : (c2041 || c2042) ? point0_ip2 : c1988 ? point0_ip2 : c1989 ? point0_ip2 : c1990 ? point0_ip2 : c1991 ? point0_ip2 : c1992 ? point0_ip2 : c1993 ? point0_ip2 : c1994 ? point0_ip2 : c1995 ? point0_ip2 : c1996 ? point0_ip2 : ((c2055 || c2091) || c2090) ? point0_ip2 : c1998 ? point0_ip2 : c1999 ? point0_ip2 : c2000 ? point0_ip2 : c2001 ? point0_ip2 : (c2199 || c2198) ? point0_ip2 : (c2002 && !c927) ? point0_ip2 : c1972 ? point0_ip2 : 'bz;
  assign point0_ip_saved4 = c2037 ? ip2 : c2038 ? point0_ip_saved2 : c2039 ? point0_ip_saved2 : c2040 ? point0_ip_saved2 : 'bz;
  assign point0_ip_saved5 = (c1971 && c889) ? point0_ip_saved2 : ((c2004 || c2005) || c2006) ? point0_ip_saved2 : c1974 ? point0_ip_saved2 : c1975 ? point0_ip_saved2 : c1976 ? point0_ip_saved2 : c1977 ? point0_ip_saved2 : c1978 ? point0_ip_saved2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? point0_ip_saved2 : (((c2019 || c2017) || c2018) || c2016) ? point0_ip_saved2 : c1981 ? point0_ip_saved2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? point0_ip_saved2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? point0_ip_saved2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? point0_ip_saved2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? point0_ip_saved2 : (((c2038 || c2040) || c2037) || c2039) ? point0_ip_saved4 : (c2041 || c2042) ? point0_ip_saved2 : c1988 ? point0_ip_saved2 : c1989 ? point0_ip_saved2 : c1990 ? point0_ip_saved2 : c1991 ? point0_ip_saved2 : c1992 ? point0_ip_saved2 : c1993 ? point0_ip_saved2 : c1994 ? point0_ip_saved2 : c1995 ? point0_ip_saved2 : c1996 ? point0_ip_saved2 : ((c2055 || c2091) || c2090) ? point0_ip_saved2 : c1998 ? point0_ip_saved2 : c1999 ? point0_ip_saved2 : c2000 ? point0_ip_saved2 : c2001 ? point0_ip_saved2 : (c2199 || c2198) ? point0_ip_saved2 : (c2002 && !c927) ? point0_ip_saved2 : c1972 ? point0_ip_saved2 : 'bz;
  assign point0_phase7 = c2037 ? 1 : c2038 ? 2 : c2039 ? 3 : c2040 ? 0 : 'bz;
  assign point0_phase8 = (c1971 && c889) ? point0_phase2 : ((c2004 || c2005) || c2006) ? point0_phase2 : c1974 ? point0_phase2 : c1975 ? point0_phase2 : c1976 ? point0_phase2 : c1977 ? point0_phase2 : c1978 ? point0_phase2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? point0_phase2 : (((c2019 || c2017) || c2018) || c2016) ? point0_phase2 : c1981 ? point0_phase2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? point0_phase2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? point0_phase2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? point0_phase2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? point0_phase2 : (((c2038 || c2040) || c2037) || c2039) ? point0_phase7 : (c2041 || c2042) ? point0_phase2 : c1988 ? point0_phase2 : c1989 ? point0_phase2 : c1990 ? point0_phase2 : c1991 ? point0_phase2 : c1992 ? point0_phase2 : c1993 ? point0_phase2 : c1994 ? point0_phase2 : c1995 ? point0_phase2 : c1996 ? point0_phase2 : ((c2055 || c2091) || c2090) ? point0_phase2 : c1998 ? point0_phase2 : c1999 ? point0_phase2 : c2000 ? point0_phase2 : c2001 ? point0_phase2 : (c2199 || c2198) ? point0_phase2 : (c2002 && !c927) ? point0_phase2 : c1972 ? point0_phase2 : 'bz;
  assign q_inl522 = (t1006_inl1_inl52 / t1006_inl2_inl52);
  assign q_inl523 = (q_inl522 * -1);
  assign q_inl524 = (q_inl522 * -1);
  assign q_inl525 = c2046 ? q_inl522 : c2047 ? q_inl523 : c2048 ? q_inl524 : (c1991 && c1096_inl52) ? q_inl522 : 'bz;
  assign r_inl522 = (t1006_inl1_inl52 % t1006_inl2_inl52);
  assign r_inl523 = (r_inl522 * -1);
  assign r_inl524 = (r_inl522 * -1);
  assign r_inl525 = c2046 ? r_inl523 : c2047 ? r_inl522 : c2048 ? r_inl524 : (c1991 && c1096_inl52) ? r_inl522 : 'bz;
  assign retro_divmod_result522[0] = array1007_inl52[0];
  assign retro_divmod_result522[1] = array1007_inl52[1];
  assign stack0_pos10 = c2124 ? stack0_pos2 : c2125 ? stack0_pos9 : c2013 ? stack0_pos2 : c2014 ? stack0_pos2 : c2015 ? stack0_pos2 : 'bz;
  assign stack0_pos11 = (stack0_pos2 - 1);
  assign stack0_pos12 = (stack0_pos2 - 1);
  assign stack0_pos13 = c2021 ? stack0_pos11 : c2022 ? stack0_pos12 : c2023 ? stack0_pos2 : c2024 ? stack0_pos2 : 'bz;
  assign stack0_pos14 = (stack0_pos2 - 1);
  assign stack0_pos15 = (stack0_pos2 - 1);
  assign stack0_pos16 = c2025 ? stack0_pos14 : c2026 ? stack0_pos15 : c2027 ? stack0_pos2 : c2028 ? stack0_pos2 : 'bz;
  assign stack0_pos17 = (stack0_pos2 - 1);
  assign stack0_pos18 = (stack0_pos2 - 1);
  assign stack0_pos19 = c2029 ? stack0_pos17 : c2030 ? stack0_pos18 : c2031 ? stack0_pos2 : c2032 ? stack0_pos2 : 'bz;
  assign stack0_pos20 = (stack0_pos2 - 1);
  assign stack0_pos21 = (stack0_pos2 - 1);
  assign stack0_pos22 = c2033 ? stack0_pos20 : c2034 ? stack0_pos21 : c2035 ? stack0_pos2 : c2036 ? stack0_pos2 : 'bz;
  assign stack0_pos23 = (stack0_pos2 - 1);
  assign stack0_pos24 = (stack0_pos2 - 1);
  assign stack0_pos25 = c2041 ? stack0_pos23 : c2042 ? stack0_pos24 : 'bz;
  assign stack0_pos26 = (stack0_pos2 - 1);
  assign stack0_pos27 = (stack0_pos2 - 1);
  assign stack0_pos28 = (stack0_pos2 - 1);
  assign stack0_pos29 = (stack0_pos2 - 1);
  assign stack0_pos30 = (stack0_pos2 - 1);
  assign stack0_pos31 = (stack0_pos2 - 1);
  assign stack0_pos32 = (stack0_pos2 - 1);
  assign stack0_pos33 = (stack0_pos2 - 1);
  assign stack0_pos34 = (stack0_pos2 - 1);
  assign stack0_pos35 = c2090 ? stack0_pos34 : c2091 ? stack0_pos2 : c2055 ? stack0_pos2 : 'bz;
  assign stack0_pos36 = (stack0_pos2 - 1);
  assign stack0_pos37 = (stack0_pos36 - 1);
  assign stack0_pos38 = (stack0_pos2 - 1);
  assign stack0_pos39 = (stack0_pos2 - 1);
  assign stack0_pos3 = (stack0_pos2 + 1);
  assign stack0_pos40 = (stack0_pos2 - 1);
  assign stack0_pos41 = c2155 ? stack0_pos38 : c2156 ? stack0_pos39 : c2152 ? stack0_pos40 : 'bz;
  assign stack0_pos42 = ((c2152 || c2155) || c2156) ? stack0_pos41 : (((c2139 || c2140) || c2120) && !c935_inl55) ? stack0_pos2 : 'bz;
  assign stack0_pos43 = (c1971 && c889) ? stack0_pos2 : ((c2004 || c2005) || c2006) ? stack0_pos4 : c1974 ? stack0_pos5 : c1975 ? stack0_pos6 : c1976 ? stack0_pos2 : c1977 ? stack0_pos7 : c1978 ? stack0_pos8 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? stack0_pos10 : (((c2019 || c2017) || c2018) || c2016) ? stack0_pos2 : c1981 ? stack0_pos2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? stack0_pos13 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? stack0_pos16 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? stack0_pos19 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? stack0_pos22 : (((c2038 || c2040) || c2037) || c2039) ? stack0_pos2 : (c2041 || c2042) ? stack0_pos25 : c1988 ? stack0_pos26 : c1989 ? stack0_pos27 : c1990 ? stack0_pos28 : c1991 ? stack0_pos2 : c1992 ? stack0_pos29 : c1993 ? stack0_pos30 : c1994 ? stack0_pos31 : c1995 ? stack0_pos32 : c1996 ? stack0_pos33 : ((c2055 || c2091) || c2090) ? stack0_pos35 : c1998 ? stack0_pos2 : c1999 ? stack0_pos2 : c2000 ? stack0_pos2 : c2001 ? stack0_pos37 : (c2199 || c2198) ? stack0_pos42 : (c2002 && !c927) ? stack0_pos2 : c1972 ? stack0_pos2 : 'bz;
  assign stack0_pos4 = c2004 ? stack0_pos2 : c2005 ? stack0_pos2 : c2006 ? stack0_pos3 : 'bz;
  assign stack0_pos5 = (stack0_pos2 + 1);
  assign stack0_pos6 = (stack0_pos2 - 1);
  assign stack0_pos7 = (stack0_pos2 - 1);
  assign stack0_pos8 = (stack0_pos2 + 1);
  assign stack0_pos9 = (stack0_pos2 - 1);
  assign stack0_second11 = c2124 ? stack0_second2 : c2125 ? stack0_second10 : c2013 ? stack0_second2 : c2014 ? stack0_second2 : c2015 ? stack0_second2 : 'bz;
  assign stack0_second14 = c2021 ? stack0_second12 : c2022 ? stack0_second13 : c2023 ? stack0_second2 : c2024 ? stack0_second2 : 'bz;
  assign stack0_second17 = c2025 ? stack0_second15 : c2026 ? stack0_second16 : c2027 ? stack0_second2 : c2028 ? stack0_second2 : 'bz;
  assign stack0_second20 = c2029 ? stack0_second18 : c2030 ? stack0_second19 : c2031 ? stack0_second2 : c2032 ? stack0_second2 : 'bz;
  assign stack0_second23 = c2033 ? stack0_second21 : c2034 ? stack0_second22 : c2035 ? stack0_second2 : c2036 ? stack0_second2 : 'bz;
  assign stack0_second26 = c2041 ? stack0_second24 : c2042 ? stack0_second25 : 'bz;
  assign stack0_second30 = retro_divmod_result522[1];
  assign stack0_second37 = c2090 ? stack0_second36 : c2091 ? stack0_second2 : c2055 ? stack0_second2 : 'bz;
  assign stack0_second43 = c2155 ? stack0_second40 : c2156 ? stack0_second41 : c2152 ? stack0_second42 : 'bz;
  assign stack0_second44 = ((c2152 || c2155) || c2156) ? stack0_second43 : (((c2139 || c2140) || c2120) && !c935_inl55) ? stack0_second2 : 'bz;
  assign stack0_second45 = (c1971 && c889) ? stack0_second2 : ((c2004 || c2005) || c2006) ? stack0_second4 : c1974 ? stack0_top2 : c1975 ? stack0_second6 : c1976 ? stack0_top2 : c1977 ? stack0_second8 : c1978 ? stack0_top2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? stack0_second11 : (((c2019 || c2017) || c2018) || c2016) ? stack0_second2 : c1981 ? stack0_second2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? stack0_second14 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? stack0_second17 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? stack0_second20 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? stack0_second23 : (((c2038 || c2040) || c2037) || c2039) ? stack0_second2 : (c2041 || c2042) ? stack0_second26 : c1988 ? stack0_second27 : c1989 ? stack0_second28 : c1990 ? stack0_second29 : c1991 ? stack0_second30 : c1992 ? stack0_second31 : c1993 ? stack0_second32 : c1994 ? stack0_second33 : c1995 ? stack0_second34 : c1996 ? stack0_second35 : ((c2055 || c2091) || c2090) ? stack0_second37 : c1998 ? stack0_second2 : c1999 ? stack0_second2 : c2000 ? stack0_second2 : c2001 ? stack0_second39 : (c2199 || c2198) ? stack0_second44 : (c2002 && !c927) ? stack0_second2 : c1972 ? stack0_second2 : 'bz;
  assign stack0_second4 = c2004 ? stack0_second2 : c2005 ? stack0_second2 : c2006 ? stack0_top2 : 'bz;
  assign stack0_top10 = (stack0_top2 - 1);
  assign stack0_top12 = c2124 ? stack0_top10 : c2125 ? stack0_second2 : c2013 ? stack0_top2 : c2014 ? stack0_top2 : c2015 ? stack0_top2 : 'bz;
  assign stack0_top15 = c2021 ? stack0_second2 : c2022 ? stack0_second2 : c2023 ? stack0_top2 : c2024 ? stack0_top2 : 'bz;
  assign stack0_top18 = c2025 ? stack0_second2 : c2026 ? stack0_second2 : c2027 ? stack0_top2 : c2028 ? stack0_top2 : 'bz;
  assign stack0_top21 = c2029 ? stack0_second2 : c2030 ? stack0_second2 : c2031 ? stack0_top2 : c2032 ? stack0_top2 : 'bz;
  assign stack0_top24 = c2033 ? stack0_second2 : c2034 ? stack0_second2 : c2035 ? stack0_top2 : c2036 ? stack0_top2 : 'bz;
  assign stack0_top26 = c2037 ? stack0_top2 : c2038 ? stack0_top2 : c2039 ? mem_data : c2040 ? stack0_top2 : 'bz;
  assign stack0_top31 = (stack0_second2 + stack0_top2);
  assign stack0_top33 = (stack0_second2 - stack0_top2);
  assign stack0_top35 = (stack0_second2 * stack0_top2);
  assign stack0_top36 = retro_divmod_result522[0];
  assign stack0_top38 = (stack0_second2 & stack0_top2);
  assign stack0_top40 = (stack0_second2 | stack0_top2);
  assign stack0_top42 = (stack0_second2 ^ stack0_top2);
  assign stack0_top44 = (stack0_second2 << stack0_top2);
  assign stack0_top46 = (stack0_second2 >>> stack0_top2);
  assign stack0_top48 = c2090 ? stack0_second2 : c2091 ? stack0_top2 : c2055 ? stack0_top2 : 'bz;
  assign stack0_top49 = (stack0_top2 + 1);
  assign stack0_top4 = c2004 ? stack0_top2 : c2005 ? stack0_top2 : c2006 ? mem_data : 'bz;
  assign stack0_top50 = (stack0_top2 - 1);
  assign stack0_top58 = ((c2152 || c2155) || c2156) ? stack0_second2 : (((c2139 || c2140) || c2120) && !c935_inl55) ? stack0_top2 : 'bz;
  assign stack0_top59 = (c1971 && c889) ? stack0_top2 : ((c2004 || c2005) || c2006) ? stack0_top4 : c1974 ? stack0_top2 : c1975 ? stack0_second2 : c1976 ? stack0_second2 : c1977 ? stack0_second2 : c1978 ? address0_top2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? stack0_top12 : (((c2019 || c2017) || c2018) || c2016) ? stack0_top2 : c1981 ? stack0_top2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? stack0_top15 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? stack0_top18 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? stack0_top21 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? stack0_top24 : (((c2038 || c2040) || c2037) || c2039) ? stack0_top26 : (c2041 || c2042) ? stack0_second2 : c1988 ? stack0_top31 : c1989 ? stack0_top33 : c1990 ? stack0_top35 : c1991 ? stack0_top36 : c1992 ? stack0_top38 : c1993 ? stack0_top40 : c1994 ? stack0_top42 : c1995 ? stack0_top44 : c1996 ? stack0_top46 : ((c2055 || c2091) || c2090) ? stack0_top48 : c1998 ? stack0_top49 : c1999 ? stack0_top50 : c2000 ? stack0_top51 : c2001 ? stack0_second38 : (c2199 || c2198) ? stack0_top58 : (c2002 && !c927) ? stack0_top2 : c1972 ? stack0_top2 : 'bz;
  assign t1006_inl1_inl52 = c1005_inl1_inl52 ? -stack0_second2 : stack0_second2;
  assign t1006_inl2_inl52 = c1005_inl2_inl52 ? -stack0_top2 : stack0_top2;
  assign t2771 = c2126 ? 0 : c2127 ? 1 : 'bz;
  assign t2774 = c2126 ? 2 : c2127 ? 0 : 'bz;
  assign t2778 = c2128 ? 0 : c2129 ? 1 : 'bz;
  assign t2781 = c2128 ? 2 : c2129 ? 0 : 'bz;
  assign t2785 = c2130 ? 0 : c2131 ? 1 : 'bz;
  assign t2788 = c2130 ? 2 : c2131 ? 0 : 'bz;
  assign t2792 = c2132 ? 0 : c2133 ? 1 : 'bz;
  assign t2795 = c2132 ? 2 : c2133 ? 0 : 'bz;
  assign t2829 = c2146 ? 1 : ((c2041 || c2042) && !c924) ? wr_flag2 : 'bz;
  assign t2830 = c2146 ? write_point0_addr4 : ((c2041 || c2042) && !c924) ? wr_mem_addr2 : 'bz;
  assign t2831 = c2146 ? write_point0_data4 : ((c2041 || c2042) && !c924) ? wr_mem_data2 : 'bz;
  assign t839_inl14 = (stack0_pos2 - 2);
  assign t839_inl15 = (address0_pos2 - 2);
  assign t839_inl16 = (stack0_pos2 - 2);
  assign t839_inl17 = (address0_pos2 - 2);
  assign t839_inl1_inl13 = (stack0_pos2 - 2);
  assign t842_inl18 = (stack0_pos6 - 2);
  assign t842_inl19 = (stack0_pos7 - 2);
  assign t842_inl1_inl35 = (stack0_pos11 - 2);
  assign t842_inl1_inl36 = (stack0_pos14 - 2);
  assign t842_inl1_inl37 = (stack0_pos17 - 2);
  assign t842_inl1_inl38 = (stack0_pos20 - 2);
  assign t842_inl1_inl40 = (stack0_pos23 - 2);
  assign t842_inl1_inl54 = (stack0_pos34 - 2);
  assign t842_inl20 = (address0_pos4 - 2);
  assign t842_inl21 = (address0_pos5 - 2);
  assign t842_inl22 = (stack0_pos26 - 2);
  assign t842_inl23 = (stack0_pos27 - 2);
  assign t842_inl24 = (stack0_pos28 - 2);
  assign t842_inl25 = (stack0_pos29 - 2);
  assign t842_inl26 = (stack0_pos30 - 2);
  assign t842_inl27 = (stack0_pos31 - 2);
  assign t842_inl28 = (stack0_pos32 - 2);
  assign t842_inl29 = (stack0_pos33 - 2);
  assign t842_inl2_inl33 = (stack0_pos9 - 2);
  assign t842_inl2_inl35 = (stack0_pos12 - 2);
  assign t842_inl2_inl36 = (stack0_pos15 - 2);
  assign t842_inl2_inl37 = (stack0_pos18 - 2);
  assign t842_inl2_inl38 = (stack0_pos21 - 2);
  assign t842_inl2_inl40 = (stack0_pos24 - 2);
  assign t842_inl2_inl54 = (address0_pos6 - 2);
  assign t842_inl2_inl55 = (stack0_pos38 - 2);
  assign t842_inl30 = (stack0_pos36 - 2);
  assign t842_inl31 = (stack0_pos37 - 2);
  assign t842_inl3_inl55 = (stack0_pos39 - 2);
  assign t842_inl4_inl55 = (stack0_pos40 - 2);
  assign wr_flag4 = (c1971 && c889) ? wr_flag2 : ((c2004 || c2005) || c2006) ? wr_flag2 : c1974 ? wr_flag2 : c1975 ? wr_flag2 : c1976 ? wr_flag2 : c1977 ? wr_flag2 : c1978 ? wr_flag2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? wr_flag2 : (((c2019 || c2017) || c2018) || c2016) ? wr_flag2 : c1981 ? wr_flag2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? wr_flag2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? wr_flag2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? wr_flag2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? wr_flag2 : (((c2038 || c2040) || c2037) || c2039) ? wr_flag2 : (c2041 || c2042) ? t2829 : c1988 ? wr_flag2 : c1989 ? wr_flag2 : c1990 ? wr_flag2 : c1991 ? wr_flag2 : c1992 ? wr_flag2 : c1993 ? wr_flag2 : c1994 ? wr_flag2 : c1995 ? wr_flag2 : c1996 ? wr_flag2 : ((c2055 || c2091) || c2090) ? wr_flag2 : c1998 ? wr_flag2 : c1999 ? wr_flag2 : c2000 ? wr_flag2 : c2001 ? wr_flag2 : (c2199 || c2198) ? wr_flag2 : (c2002 && !c927) ? wr_flag2 : c1972 ? wr_flag2 : 'bz;
  assign wr_flag6 = c2200 ? 0 : (c886 && !c920) ? wr_flag4 : 'bz;
  assign wr_mem_addr4 = (c1971 && c889) ? wr_mem_addr2 : ((c2004 || c2005) || c2006) ? wr_mem_addr2 : c1974 ? wr_mem_addr2 : c1975 ? wr_mem_addr2 : c1976 ? wr_mem_addr2 : c1977 ? wr_mem_addr2 : c1978 ? wr_mem_addr2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? wr_mem_addr2 : (((c2019 || c2017) || c2018) || c2016) ? wr_mem_addr2 : c1981 ? wr_mem_addr2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? wr_mem_addr2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? wr_mem_addr2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? wr_mem_addr2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? wr_mem_addr2 : (((c2038 || c2040) || c2037) || c2039) ? wr_mem_addr2 : (c2041 || c2042) ? t2830 : c1988 ? wr_mem_addr2 : c1989 ? wr_mem_addr2 : c1990 ? wr_mem_addr2 : c1991 ? wr_mem_addr2 : c1992 ? wr_mem_addr2 : c1993 ? wr_mem_addr2 : c1994 ? wr_mem_addr2 : c1995 ? wr_mem_addr2 : c1996 ? wr_mem_addr2 : ((c2055 || c2091) || c2090) ? wr_mem_addr2 : c1998 ? wr_mem_addr2 : c1999 ? wr_mem_addr2 : c2000 ? wr_mem_addr2 : c2001 ? wr_mem_addr2 : (c2199 || c2198) ? wr_mem_addr2 : (c2002 && !c927) ? wr_mem_addr2 : c1972 ? wr_mem_addr2 : 'bz;
  assign wr_mem_data4 = (c1971 && c889) ? wr_mem_data2 : ((c2004 || c2005) || c2006) ? wr_mem_data2 : c1974 ? wr_mem_data2 : c1975 ? wr_mem_data2 : c1976 ? wr_mem_data2 : c1977 ? wr_mem_data2 : c1978 ? wr_mem_data2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? wr_mem_data2 : (((c2019 || c2017) || c2018) || c2016) ? wr_mem_data2 : c1981 ? wr_mem_data2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? wr_mem_data2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? wr_mem_data2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? wr_mem_data2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? wr_mem_data2 : (((c2038 || c2040) || c2037) || c2039) ? wr_mem_data2 : (c2041 || c2042) ? t2831 : c1988 ? wr_mem_data2 : c1989 ? wr_mem_data2 : c1990 ? wr_mem_data2 : c1991 ? wr_mem_data2 : c1992 ? wr_mem_data2 : c1993 ? wr_mem_data2 : c1994 ? wr_mem_data2 : c1995 ? wr_mem_data2 : c1996 ? wr_mem_data2 : ((c2055 || c2091) || c2090) ? wr_mem_data2 : c1998 ? wr_mem_data2 : c1999 ? wr_mem_data2 : c2000 ? wr_mem_data2 : c2001 ? wr_mem_data2 : (c2199 || c2198) ? wr_mem_data2 : (c2002 && !c927) ? wr_mem_data2 : c1972 ? wr_mem_data2 : 'bz;
  assign write_point0_addr4 = c2041 ? stack0_top2 : c2042 ? write_point0_addr2 : 'bz;
  assign write_point0_addr5 = (c1971 && c889) ? write_point0_addr2 : ((c2004 || c2005) || c2006) ? write_point0_addr2 : c1974 ? write_point0_addr2 : c1975 ? write_point0_addr2 : c1976 ? write_point0_addr2 : c1977 ? write_point0_addr2 : c1978 ? write_point0_addr2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? write_point0_addr2 : (((c2019 || c2017) || c2018) || c2016) ? write_point0_addr2 : c1981 ? write_point0_addr2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? write_point0_addr2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? write_point0_addr2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? write_point0_addr2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? write_point0_addr2 : (((c2038 || c2040) || c2037) || c2039) ? write_point0_addr2 : (c2041 || c2042) ? write_point0_addr4 : c1988 ? write_point0_addr2 : c1989 ? write_point0_addr2 : c1990 ? write_point0_addr2 : c1991 ? write_point0_addr2 : c1992 ? write_point0_addr2 : c1993 ? write_point0_addr2 : c1994 ? write_point0_addr2 : c1995 ? write_point0_addr2 : c1996 ? write_point0_addr2 : ((c2055 || c2091) || c2090) ? write_point0_addr2 : c1998 ? write_point0_addr2 : c1999 ? write_point0_addr2 : c2000 ? write_point0_addr2 : c2001 ? write_point0_addr2 : (c2199 || c2198) ? write_point0_addr2 : (c2002 && !c927) ? write_point0_addr2 : c1972 ? write_point0_addr2 : 'bz;
  assign write_point0_data4 = c2041 ? write_point0_data2 : c2042 ? stack0_top2 : 'bz;
  assign write_point0_data5 = (c1971 && c889) ? write_point0_data2 : ((c2004 || c2005) || c2006) ? write_point0_data2 : c1974 ? write_point0_data2 : c1975 ? write_point0_data2 : c1976 ? write_point0_data2 : c1977 ? write_point0_data2 : c1978 ? write_point0_data2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? write_point0_data2 : (((c2019 || c2017) || c2018) || c2016) ? write_point0_data2 : c1981 ? write_point0_data2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? write_point0_data2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? write_point0_data2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? write_point0_data2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? write_point0_data2 : (((c2038 || c2040) || c2037) || c2039) ? write_point0_data2 : (c2041 || c2042) ? write_point0_data4 : c1988 ? write_point0_data2 : c1989 ? write_point0_data2 : c1990 ? write_point0_data2 : c1991 ? write_point0_data2 : c1992 ? write_point0_data2 : c1993 ? write_point0_data2 : c1994 ? write_point0_data2 : c1995 ? write_point0_data2 : c1996 ? write_point0_data2 : ((c2055 || c2091) || c2090) ? write_point0_data2 : c1998 ? write_point0_data2 : c1999 ? write_point0_data2 : c2000 ? write_point0_data2 : c2001 ? write_point0_data2 : (c2199 || c2198) ? write_point0_data2 : (c2002 && !c927) ? write_point0_data2 : c1972 ? write_point0_data2 : 'bz;
  assign write_point0_ip4 = c2041 ? ip2 : c2042 ? write_point0_ip2 : 'bz;
  assign write_point0_ip5 = (c1971 && c889) ? write_point0_ip2 : ((c2004 || c2005) || c2006) ? write_point0_ip2 : c1974 ? write_point0_ip2 : c1975 ? write_point0_ip2 : c1976 ? write_point0_ip2 : c1977 ? write_point0_ip2 : c1978 ? write_point0_ip2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? write_point0_ip2 : (((c2019 || c2017) || c2018) || c2016) ? write_point0_ip2 : c1981 ? write_point0_ip2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? write_point0_ip2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? write_point0_ip2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? write_point0_ip2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? write_point0_ip2 : (((c2038 || c2040) || c2037) || c2039) ? write_point0_ip2 : (c2041 || c2042) ? write_point0_ip4 : c1988 ? write_point0_ip2 : c1989 ? write_point0_ip2 : c1990 ? write_point0_ip2 : c1991 ? write_point0_ip2 : c1992 ? write_point0_ip2 : c1993 ? write_point0_ip2 : c1994 ? write_point0_ip2 : c1995 ? write_point0_ip2 : c1996 ? write_point0_ip2 : ((c2055 || c2091) || c2090) ? write_point0_ip2 : c1998 ? write_point0_ip2 : c1999 ? write_point0_ip2 : c2000 ? write_point0_ip2 : c2001 ? write_point0_ip2 : (c2199 || c2198) ? write_point0_ip2 : (c2002 && !c927) ? write_point0_ip2 : c1972 ? write_point0_ip2 : 'bz;
  assign write_point0_phase5 = c2041 ? 1 : c2042 ? 0 : 'bz;
  assign write_point0_phase6 = (c1971 && c889) ? write_point0_phase2 : ((c2004 || c2005) || c2006) ? write_point0_phase2 : c1974 ? write_point0_phase2 : c1975 ? write_point0_phase2 : c1976 ? write_point0_phase2 : c1977 ? write_point0_phase2 : c1978 ? write_point0_phase2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? write_point0_phase2 : (((c2019 || c2017) || c2018) || c2016) ? write_point0_phase2 : c1981 ? write_point0_phase2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? write_point0_phase2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? write_point0_phase2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? write_point0_phase2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? write_point0_phase2 : (((c2038 || c2040) || c2037) || c2039) ? write_point0_phase2 : (c2041 || c2042) ? write_point0_phase5 : c1988 ? write_point0_phase2 : c1989 ? write_point0_phase2 : c1990 ? write_point0_phase2 : c1991 ? write_point0_phase2 : c1992 ? write_point0_phase2 : c1993 ? write_point0_phase2 : c1994 ? write_point0_phase2 : c1995 ? write_point0_phase2 : c1996 ? write_point0_phase2 : ((c2055 || c2091) || c2090) ? write_point0_phase2 : c1998 ? write_point0_phase2 : c1999 ? write_point0_phase2 : c2000 ? write_point0_phase2 : c2001 ? write_point0_phase2 : (c2199 || c2198) ? write_point0_phase2 : (c2002 && !c927) ? write_point0_phase2 : c1972 ? write_point0_phase2 : 'bz;
  assign zero_pop_return0_ip5 = c2090 ? address0_top2 : c2091 ? ip2 : c2055 ? zero_pop_return0_ip2 : 'bz;
  assign zero_pop_return0_ip6 = (c1971 && c889) ? zero_pop_return0_ip2 : ((c2004 || c2005) || c2006) ? zero_pop_return0_ip2 : c1974 ? zero_pop_return0_ip2 : c1975 ? zero_pop_return0_ip2 : c1976 ? zero_pop_return0_ip2 : c1977 ? zero_pop_return0_ip2 : c1978 ? zero_pop_return0_ip2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? zero_pop_return0_ip2 : (((c2019 || c2017) || c2018) || c2016) ? zero_pop_return0_ip2 : c1981 ? zero_pop_return0_ip2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? zero_pop_return0_ip2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? zero_pop_return0_ip2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? zero_pop_return0_ip2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? zero_pop_return0_ip2 : (((c2038 || c2040) || c2037) || c2039) ? zero_pop_return0_ip2 : (c2041 || c2042) ? zero_pop_return0_ip2 : c1988 ? zero_pop_return0_ip2 : c1989 ? zero_pop_return0_ip2 : c1990 ? zero_pop_return0_ip2 : c1991 ? zero_pop_return0_ip2 : c1992 ? zero_pop_return0_ip2 : c1993 ? zero_pop_return0_ip2 : c1994 ? zero_pop_return0_ip2 : c1995 ? zero_pop_return0_ip2 : c1996 ? zero_pop_return0_ip2 : ((c2055 || c2091) || c2090) ? zero_pop_return0_ip5 : c1998 ? zero_pop_return0_ip2 : c1999 ? zero_pop_return0_ip2 : c2000 ? zero_pop_return0_ip2 : c2001 ? zero_pop_return0_ip2 : (c2199 || c2198) ? zero_pop_return0_ip2 : (c2002 && !c927) ? zero_pop_return0_ip2 : c1972 ? zero_pop_return0_ip2 : 'bz;
  assign zero_pop_return0_phase5 = c2090 ? 1 : c2091 ? zero_pop_return0_phase2 : c2055 ? 0 : 'bz;
  assign zero_pop_return0_phase6 = (c1971 && c889) ? zero_pop_return0_phase2 : ((c2004 || c2005) || c2006) ? zero_pop_return0_phase2 : c1974 ? zero_pop_return0_phase2 : c1975 ? zero_pop_return0_phase2 : c1976 ? zero_pop_return0_phase2 : c1977 ? zero_pop_return0_phase2 : c1978 ? zero_pop_return0_phase2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? zero_pop_return0_phase2 : (((c2019 || c2017) || c2018) || c2016) ? zero_pop_return0_phase2 : c1981 ? zero_pop_return0_phase2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? zero_pop_return0_phase2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? zero_pop_return0_phase2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? zero_pop_return0_phase2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? zero_pop_return0_phase2 : (((c2038 || c2040) || c2037) || c2039) ? zero_pop_return0_phase2 : (c2041 || c2042) ? zero_pop_return0_phase2 : c1988 ? zero_pop_return0_phase2 : c1989 ? zero_pop_return0_phase2 : c1990 ? zero_pop_return0_phase2 : c1991 ? zero_pop_return0_phase2 : c1992 ? zero_pop_return0_phase2 : c1993 ? zero_pop_return0_phase2 : c1994 ? zero_pop_return0_phase2 : c1995 ? zero_pop_return0_phase2 : c1996 ? zero_pop_return0_phase2 : ((c2055 || c2091) || c2090) ? zero_pop_return0_phase5 : c1998 ? zero_pop_return0_phase2 : c1999 ? zero_pop_return0_phase2 : c2000 ? zero_pop_return0_phase2 : c2001 ? zero_pop_return0_phase2 : (c2199 || c2198) ? zero_pop_return0_phase2 : (c2002 && !c927) ? zero_pop_return0_phase2 : c1972 ? zero_pop_return0_phase2 : 'bz;
  //combinations: array1008
  assign _stack_len = array1008_ram_len;
  assign _stack_q = array1008_ram_q;
  assign array1008_ram_addr = _stack_addr;
  assign array1008_ram_d = _stack_d;
  assign array1008_ram_we = _stack_we;
  //combinations: array1009
  assign _address_len = array1009_ram_len;
  assign _address_q = array1009_ram_q;
  assign array1009_ram_addr = _address_addr;
  assign array1009_ram_d = _address_d;
  assign array1009_ram_we = _address_we;
  //combinations: in_io_ports
  assign io_ports_len = retro_main_in_io_ports_len;
  assign io_ports_q = retro_main_in_io_ports_q;
  assign retro_main_in_io_ports_addr = io_ports_addr;
  assign retro_main_in_io_ports_d = io_ports_d;
  assign retro_main_in_io_ports_req = io_ports_req;
  assign retro_main_in_io_ports_we = io_ports_we;
  //combinations: in_memory
  assign memory_len = retro_main_in_memory_len;
  assign memory_q = retro_main_in_memory_q;
  assign retro_main_in_memory_addr = memory_addr;
  assign retro_main_in_memory_d = memory_d;
  assign retro_main_in_memory_req = memory_req;
  assign retro_main_in_memory_we = memory_we;
  //sub modules
  //array1008 instance
  BidirectionalSinglePortRam#(
    .DATA_WIDTH(32),
    .ADDR_WIDTH(8),
    .RAM_LENGTH(128)
    )
    array1008(
      .clk(clk),
      .rst(rst),
      .ram_addr(array1008_ram_addr),
      .ram_d(array1008_ram_d),
      .ram_we(array1008_ram_we),
      .ram_q(array1008_ram_q),
      .ram_len(array1008_ram_len)
    );
  //array1009 instance
  BidirectionalSinglePortRam#(
    .DATA_WIDTH(32),
    .ADDR_WIDTH(11),
    .RAM_LENGTH(1024)
    )
    array1009(
      .clk(clk),
      .rst(rst),
      .ram_addr(array1009_ram_addr),
      .ram_d(array1009_ram_d),
      .ram_we(array1009_ram_we),
      .ram_q(array1009_ram_q),
      .ram_len(array1009_ram_len)
    );
  
  
  always @(posedge clk) begin
    if (rst) begin
      _address_addr <= 0;
      _address_d <= 0;
      _address_req <= 0;
      _address_we <= 0;
      _stack_addr <= 0;
      _stack_d <= 0;
      _stack_req <= 0;
      _stack_we <= 0;
      address0_pos2 <= 0;
      address0_second2 <= 0;
      address0_second4 <= 0;
      address0_second5 <= 0;
      address0_second6 <= 0;
      address0_top2 <= 0;
      done_flag2 <= 0;
      exec_result336 <= 0;
      io_ports_addr <= 0;
      io_ports_d <= 0;
      io_ports_req <= 0;
      io_ports_we <= 0;
      ip2 <= 0;
      jump0_ip2 <= 0;
      jump0_phase2 <= 0;
      jump_eq0_a2 <= 0;
      jump_eq0_ip2 <= 0;
      jump_eq0_phase2 <= 0;
      jump_ge0_a2 <= 0;
      jump_ge0_ip2 <= 0;
      jump_ge0_phase2 <= 0;
      jump_le0_a2 <= 0;
      jump_le0_ip2 <= 0;
      jump_le0_phase2 <= 0;
      jump_ne0_a2 <= 0;
      jump_ne0_ip2 <= 0;
      jump_ne0_phase2 <= 0;
      lit0_ip2 <= 0;
      lit0_phase2 <= 0;
      loop0_ip2 <= 0;
      loop0_phase2 <= 0;
      mem_data <= 0;
      memory_addr <= 0;
      memory_d <= 0;
      memory_req <= 0;
      memory_we <= 0;
      opcode2 <= 0;
      point0_ip2 <= 0;
      point0_ip_saved2 <= 0;
      point0_phase2 <= 0;
      stack0_pos2 <= 0;
      stack0_second10 <= 0;
      stack0_second12 <= 0;
      stack0_second13 <= 0;
      stack0_second15 <= 0;
      stack0_second16 <= 0;
      stack0_second18 <= 0;
      stack0_second19 <= 0;
      stack0_second21 <= 0;
      stack0_second22 <= 0;
      stack0_second24 <= 0;
      stack0_second25 <= 0;
      stack0_second27 <= 0;
      stack0_second28 <= 0;
      stack0_second29 <= 0;
      stack0_second2 <= 0;
      stack0_second31 <= 0;
      stack0_second32 <= 0;
      stack0_second33 <= 0;
      stack0_second34 <= 0;
      stack0_second35 <= 0;
      stack0_second36 <= 0;
      stack0_second38 <= 0;
      stack0_second39 <= 0;
      stack0_second40 <= 0;
      stack0_second41 <= 0;
      stack0_second42 <= 0;
      stack0_second6 <= 0;
      stack0_second8 <= 0;
      stack0_top2 <= 0;
      stack0_top51 <= 0;
      t11 <= 0;
      t926 <= 0;
      t928 <= 0;
      t929_inl55 <= 0;
      t932_inl55 <= 0;
      t934_inl55 <= 0;
      t941_inl55 <= 0;
      t943_inl55 <= 0;
      t945_inl55 <= 0;
      t947_inl55 <= 0;
      t949_inl55 <= 0;
      t951_inl55 <= 0;
      t953_inl55 <= 0;
      t955_inl55 <= 0;
      t957_inl55 <= 0;
      t959_inl55 <= 0;
      t961_inl55 <= 0;
      t963_inl55 <= 0;
      t965_inl55 <= 0;
      t967_inl55 <= 0;
      t969_inl55 <= 0;
      t971_inl55 <= 0;
      t973_inl55 <= 0;
      t975_inl55 <= 0;
      t977_inl55 <= 0;
      t979_inl55 <= 0;
      t981_inl55 <= 0;
      t983_inl55 <= 0;
      t985_inl55 <= 0;
      t987_inl55 <= 0;
      t989_inl55 <= 0;
      t991_inl55 <= 0;
      wr_flag2 <= 0;
      wr_mem_addr2 <= 0;
      wr_mem_data2 <= 0;
      write_point0_addr2 <= 0;
      write_point0_data2 <= 0;
      write_point0_ip2 <= 0;
      write_point0_phase2 <= 0;
      zero_pop_return0_ip2 <= 0;
      zero_pop_return0_phase2 <= 0;
      retro_main_state <= retro_main_b1_INIT;
    end else begin //if (rst)
      case(retro_main_state)
      retro_main_b1_INIT: begin
        retro_main_valid <= 0;
        if (retro_main_ready == 1) begin
          _address_addr <= 0;
          _address_we <= 1;
          _address_req <= 1;
          _address_d <= 0;
          _stack_addr <= 0;
          _stack_we <= 1;
          _stack_req <= 1;
          _stack_d <= 0;
          array1010[0] <= 0;
          array1010[1] <= 0;
          array1010[2] <= 0;
          array1010[3] <= 0;
          array1010[4] <= 0;
          array1010[5] <= 0;
          array1010[6] <= 0;
          array1010[7] <= 0;
          array1010[8] <= 0;
          array1010[9] <= 0;
          array1010[10] <= 0;
          array1010[11] <= 0;
          address0_pos2 <= 0;
          address0_second2 <= 0;
          address0_top2 <= 0;
          done_flag2 <= 1;
          ip2 <= 0;
          jump0_ip2 <= 0;
          jump0_phase2 <= 0;
          jump_eq0_a2 <= 0;
          jump_eq0_ip2 <= 0;
          jump_eq0_phase2 <= 0;
          jump_ge0_a2 <= 0;
          jump_ge0_ip2 <= 0;
          jump_ge0_phase2 <= 0;
          jump_le0_a2 <= 0;
          jump_le0_ip2 <= 0;
          jump_le0_phase2 <= 0;
          jump_ne0_a2 <= 0;
          jump_ne0_ip2 <= 0;
          jump_ne0_phase2 <= 0;
          lit0_ip2 <= 0;
          lit0_phase2 <= 0;
          loop0_ip2 <= 0;
          loop0_phase2 <= 0;
          opcode2 <= 0;
          point0_ip2 <= 0;
          point0_ip_saved2 <= 0;
          point0_phase2 <= 0;
          stack0_pos2 <= 0;
          stack0_second2 <= 0;
          stack0_top2 <= 0;
          wr_flag2 <= 0;
          wr_mem_addr2 <= 0;
          wr_mem_data2 <= 0;
          write_point0_addr2 <= 0;
          write_point0_data2 <= 0;
          write_point0_ip2 <= 0;
          write_point0_phase2 <= 0;
          zero_pop_return0_ip2 <= 0;
          zero_pop_return0_phase2 <= 0;
          retro_main_state <= retro_main_b1_S1;
        end
      end
      retro_main_b1_S1: begin
        _address_addr <= 1;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 1;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S2;
      end
      retro_main_b1_S2: begin
        _address_addr <= 2;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 2;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S3;
      end
      retro_main_b1_S3: begin
        _address_addr <= 3;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 3;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S4;
      end
      retro_main_b1_S4: begin
        _address_addr <= 4;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 4;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S5;
      end
      retro_main_b1_S5: begin
        _address_addr <= 5;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 5;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S6;
      end
      retro_main_b1_S6: begin
        _address_addr <= 6;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 6;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S7;
      end
      retro_main_b1_S7: begin
        _address_addr <= 7;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 7;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S8;
      end
      retro_main_b1_S8: begin
        _address_addr <= 8;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 8;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S9;
      end
      retro_main_b1_S9: begin
        _address_addr <= 9;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 9;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S10;
      end
      retro_main_b1_S10: begin
        _address_addr <= 10;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 10;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S11;
      end
      retro_main_b1_S11: begin
        _address_addr <= 11;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 11;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S12;
      end
      retro_main_b1_S12: begin
        _address_addr <= 12;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 12;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S13;
      end
      retro_main_b1_S13: begin
        _address_addr <= 13;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 13;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S14;
      end
      retro_main_b1_S14: begin
        _address_addr <= 14;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 14;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S15;
      end
      retro_main_b1_S15: begin
        _address_addr <= 15;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 15;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S16;
      end
      retro_main_b1_S16: begin
        _address_addr <= 16;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 16;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S17;
      end
      retro_main_b1_S17: begin
        _address_addr <= 17;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 17;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S18;
      end
      retro_main_b1_S18: begin
        _address_addr <= 18;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 18;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S19;
      end
      retro_main_b1_S19: begin
        _address_addr <= 19;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 19;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S20;
      end
      retro_main_b1_S20: begin
        _address_addr <= 20;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 20;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S21;
      end
      retro_main_b1_S21: begin
        _address_addr <= 21;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 21;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S22;
      end
      retro_main_b1_S22: begin
        _address_addr <= 22;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 22;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S23;
      end
      retro_main_b1_S23: begin
        _address_addr <= 23;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 23;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S24;
      end
      retro_main_b1_S24: begin
        _address_addr <= 24;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 24;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S25;
      end
      retro_main_b1_S25: begin
        _address_addr <= 25;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 25;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S26;
      end
      retro_main_b1_S26: begin
        _address_addr <= 26;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 26;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S27;
      end
      retro_main_b1_S27: begin
        _address_addr <= 27;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 27;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S28;
      end
      retro_main_b1_S28: begin
        _address_addr <= 28;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 28;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S29;
      end
      retro_main_b1_S29: begin
        _address_addr <= 29;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 29;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S30;
      end
      retro_main_b1_S30: begin
        _address_addr <= 30;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 30;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S31;
      end
      retro_main_b1_S31: begin
        _address_addr <= 31;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 31;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S32;
      end
      retro_main_b1_S32: begin
        _address_addr <= 32;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 32;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S33;
      end
      retro_main_b1_S33: begin
        _address_addr <= 33;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 33;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S34;
      end
      retro_main_b1_S34: begin
        _address_addr <= 34;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 34;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S35;
      end
      retro_main_b1_S35: begin
        _address_addr <= 35;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 35;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S36;
      end
      retro_main_b1_S36: begin
        _address_addr <= 36;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 36;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S37;
      end
      retro_main_b1_S37: begin
        _address_addr <= 37;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 37;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S38;
      end
      retro_main_b1_S38: begin
        _address_addr <= 38;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 38;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S39;
      end
      retro_main_b1_S39: begin
        _address_addr <= 39;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 39;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S40;
      end
      retro_main_b1_S40: begin
        _address_addr <= 40;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 40;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S41;
      end
      retro_main_b1_S41: begin
        _address_addr <= 41;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 41;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S42;
      end
      retro_main_b1_S42: begin
        _address_addr <= 42;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 42;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S43;
      end
      retro_main_b1_S43: begin
        _address_addr <= 43;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 43;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S44;
      end
      retro_main_b1_S44: begin
        _address_addr <= 44;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 44;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S45;
      end
      retro_main_b1_S45: begin
        _address_addr <= 45;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 45;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S46;
      end
      retro_main_b1_S46: begin
        _address_addr <= 46;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 46;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S47;
      end
      retro_main_b1_S47: begin
        _address_addr <= 47;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 47;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S48;
      end
      retro_main_b1_S48: begin
        _address_addr <= 48;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 48;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S49;
      end
      retro_main_b1_S49: begin
        _address_addr <= 49;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 49;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S50;
      end
      retro_main_b1_S50: begin
        _address_addr <= 50;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 50;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S51;
      end
      retro_main_b1_S51: begin
        _address_addr <= 51;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 51;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S52;
      end
      retro_main_b1_S52: begin
        _address_addr <= 52;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 52;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S53;
      end
      retro_main_b1_S53: begin
        _address_addr <= 53;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 53;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S54;
      end
      retro_main_b1_S54: begin
        _address_addr <= 54;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 54;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S55;
      end
      retro_main_b1_S55: begin
        _address_addr <= 55;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 55;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S56;
      end
      retro_main_b1_S56: begin
        _address_addr <= 56;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 56;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S57;
      end
      retro_main_b1_S57: begin
        _address_addr <= 57;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 57;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S58;
      end
      retro_main_b1_S58: begin
        _address_addr <= 58;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 58;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S59;
      end
      retro_main_b1_S59: begin
        _address_addr <= 59;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 59;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S60;
      end
      retro_main_b1_S60: begin
        _address_addr <= 60;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 60;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S61;
      end
      retro_main_b1_S61: begin
        _address_addr <= 61;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 61;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S62;
      end
      retro_main_b1_S62: begin
        _address_addr <= 62;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 62;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S63;
      end
      retro_main_b1_S63: begin
        _address_addr <= 63;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 63;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S64;
      end
      retro_main_b1_S64: begin
        _address_addr <= 64;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 64;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S65;
      end
      retro_main_b1_S65: begin
        _address_addr <= 65;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 65;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S66;
      end
      retro_main_b1_S66: begin
        _address_addr <= 66;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 66;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S67;
      end
      retro_main_b1_S67: begin
        _address_addr <= 67;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 67;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S68;
      end
      retro_main_b1_S68: begin
        _address_addr <= 68;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 68;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S69;
      end
      retro_main_b1_S69: begin
        _address_addr <= 69;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 69;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S70;
      end
      retro_main_b1_S70: begin
        _address_addr <= 70;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 70;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S71;
      end
      retro_main_b1_S71: begin
        _address_addr <= 71;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 71;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S72;
      end
      retro_main_b1_S72: begin
        _address_addr <= 72;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 72;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S73;
      end
      retro_main_b1_S73: begin
        _address_addr <= 73;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 73;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S74;
      end
      retro_main_b1_S74: begin
        _address_addr <= 74;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 74;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S75;
      end
      retro_main_b1_S75: begin
        _address_addr <= 75;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 75;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S76;
      end
      retro_main_b1_S76: begin
        _address_addr <= 76;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 76;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S77;
      end
      retro_main_b1_S77: begin
        _address_addr <= 77;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 77;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S78;
      end
      retro_main_b1_S78: begin
        _address_addr <= 78;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 78;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S79;
      end
      retro_main_b1_S79: begin
        _address_addr <= 79;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 79;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S80;
      end
      retro_main_b1_S80: begin
        _address_addr <= 80;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 80;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S81;
      end
      retro_main_b1_S81: begin
        _address_addr <= 81;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 81;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S82;
      end
      retro_main_b1_S82: begin
        _address_addr <= 82;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 82;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S83;
      end
      retro_main_b1_S83: begin
        _address_addr <= 83;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 83;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S84;
      end
      retro_main_b1_S84: begin
        _address_addr <= 84;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 84;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S85;
      end
      retro_main_b1_S85: begin
        _address_addr <= 85;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 85;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S86;
      end
      retro_main_b1_S86: begin
        _address_addr <= 86;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 86;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S87;
      end
      retro_main_b1_S87: begin
        _address_addr <= 87;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 87;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S88;
      end
      retro_main_b1_S88: begin
        _address_addr <= 88;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 88;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S89;
      end
      retro_main_b1_S89: begin
        _address_addr <= 89;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 89;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S90;
      end
      retro_main_b1_S90: begin
        _address_addr <= 90;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 90;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S91;
      end
      retro_main_b1_S91: begin
        _address_addr <= 91;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 91;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S92;
      end
      retro_main_b1_S92: begin
        _address_addr <= 92;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 92;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S93;
      end
      retro_main_b1_S93: begin
        _address_addr <= 93;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 93;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S94;
      end
      retro_main_b1_S94: begin
        _address_addr <= 94;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 94;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S95;
      end
      retro_main_b1_S95: begin
        _address_addr <= 95;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 95;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S96;
      end
      retro_main_b1_S96: begin
        _address_addr <= 96;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 96;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S97;
      end
      retro_main_b1_S97: begin
        _address_addr <= 97;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 97;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S98;
      end
      retro_main_b1_S98: begin
        _address_addr <= 98;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 98;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S99;
      end
      retro_main_b1_S99: begin
        _address_addr <= 99;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 99;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S100;
      end
      retro_main_b1_S100: begin
        _address_addr <= 100;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 100;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S101;
      end
      retro_main_b1_S101: begin
        _address_addr <= 101;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 101;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S102;
      end
      retro_main_b1_S102: begin
        _address_addr <= 102;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 102;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S103;
      end
      retro_main_b1_S103: begin
        _address_addr <= 103;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 103;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S104;
      end
      retro_main_b1_S104: begin
        _address_addr <= 104;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 104;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S105;
      end
      retro_main_b1_S105: begin
        _address_addr <= 105;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 105;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S106;
      end
      retro_main_b1_S106: begin
        _address_addr <= 106;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 106;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S107;
      end
      retro_main_b1_S107: begin
        _address_addr <= 107;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 107;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S108;
      end
      retro_main_b1_S108: begin
        _address_addr <= 108;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 108;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S109;
      end
      retro_main_b1_S109: begin
        _address_addr <= 109;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 109;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S110;
      end
      retro_main_b1_S110: begin
        _address_addr <= 110;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 110;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S111;
      end
      retro_main_b1_S111: begin
        _address_addr <= 111;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 111;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S112;
      end
      retro_main_b1_S112: begin
        _address_addr <= 112;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 112;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S113;
      end
      retro_main_b1_S113: begin
        _address_addr <= 113;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 113;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S114;
      end
      retro_main_b1_S114: begin
        _address_addr <= 114;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 114;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S115;
      end
      retro_main_b1_S115: begin
        _address_addr <= 115;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 115;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S116;
      end
      retro_main_b1_S116: begin
        _address_addr <= 116;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 116;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S117;
      end
      retro_main_b1_S117: begin
        _address_addr <= 117;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 117;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S118;
      end
      retro_main_b1_S118: begin
        _address_addr <= 118;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 118;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S119;
      end
      retro_main_b1_S119: begin
        _address_addr <= 119;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 119;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S120;
      end
      retro_main_b1_S120: begin
        _address_addr <= 120;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 120;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S121;
      end
      retro_main_b1_S121: begin
        _address_addr <= 121;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 121;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S122;
      end
      retro_main_b1_S122: begin
        _address_addr <= 122;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 122;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S123;
      end
      retro_main_b1_S123: begin
        _address_addr <= 123;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 123;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S124;
      end
      retro_main_b1_S124: begin
        _address_addr <= 124;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 124;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S125;
      end
      retro_main_b1_S125: begin
        _address_addr <= 125;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 125;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S126;
      end
      retro_main_b1_S126: begin
        _address_addr <= 126;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 126;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S127;
      end
      retro_main_b1_S127: begin
        _address_addr <= 127;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 127;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S128;
      end
      retro_main_b1_S128: begin
        _address_addr <= 128;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_req <= 0;
        retro_main_state <= retro_main_b1_S129;
      end
      retro_main_b1_S129: begin
        _address_addr <= 129;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S130;
      end
      retro_main_b1_S130: begin
        _address_addr <= 130;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S131;
      end
      retro_main_b1_S131: begin
        _address_addr <= 131;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S132;
      end
      retro_main_b1_S132: begin
        _address_addr <= 132;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S133;
      end
      retro_main_b1_S133: begin
        _address_addr <= 133;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S134;
      end
      retro_main_b1_S134: begin
        _address_addr <= 134;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S135;
      end
      retro_main_b1_S135: begin
        _address_addr <= 135;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S136;
      end
      retro_main_b1_S136: begin
        _address_addr <= 136;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S137;
      end
      retro_main_b1_S137: begin
        _address_addr <= 137;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S138;
      end
      retro_main_b1_S138: begin
        _address_addr <= 138;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S139;
      end
      retro_main_b1_S139: begin
        _address_addr <= 139;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S140;
      end
      retro_main_b1_S140: begin
        _address_addr <= 140;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S141;
      end
      retro_main_b1_S141: begin
        _address_addr <= 141;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S142;
      end
      retro_main_b1_S142: begin
        _address_addr <= 142;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S143;
      end
      retro_main_b1_S143: begin
        _address_addr <= 143;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S144;
      end
      retro_main_b1_S144: begin
        _address_addr <= 144;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S145;
      end
      retro_main_b1_S145: begin
        _address_addr <= 145;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S146;
      end
      retro_main_b1_S146: begin
        _address_addr <= 146;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S147;
      end
      retro_main_b1_S147: begin
        _address_addr <= 147;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S148;
      end
      retro_main_b1_S148: begin
        _address_addr <= 148;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S149;
      end
      retro_main_b1_S149: begin
        _address_addr <= 149;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S150;
      end
      retro_main_b1_S150: begin
        _address_addr <= 150;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S151;
      end
      retro_main_b1_S151: begin
        _address_addr <= 151;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S152;
      end
      retro_main_b1_S152: begin
        _address_addr <= 152;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S153;
      end
      retro_main_b1_S153: begin
        _address_addr <= 153;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S154;
      end
      retro_main_b1_S154: begin
        _address_addr <= 154;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S155;
      end
      retro_main_b1_S155: begin
        _address_addr <= 155;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S156;
      end
      retro_main_b1_S156: begin
        _address_addr <= 156;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S157;
      end
      retro_main_b1_S157: begin
        _address_addr <= 157;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S158;
      end
      retro_main_b1_S158: begin
        _address_addr <= 158;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S159;
      end
      retro_main_b1_S159: begin
        _address_addr <= 159;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S160;
      end
      retro_main_b1_S160: begin
        _address_addr <= 160;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S161;
      end
      retro_main_b1_S161: begin
        _address_addr <= 161;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S162;
      end
      retro_main_b1_S162: begin
        _address_addr <= 162;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S163;
      end
      retro_main_b1_S163: begin
        _address_addr <= 163;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S164;
      end
      retro_main_b1_S164: begin
        _address_addr <= 164;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S165;
      end
      retro_main_b1_S165: begin
        _address_addr <= 165;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S166;
      end
      retro_main_b1_S166: begin
        _address_addr <= 166;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S167;
      end
      retro_main_b1_S167: begin
        _address_addr <= 167;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S168;
      end
      retro_main_b1_S168: begin
        _address_addr <= 168;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S169;
      end
      retro_main_b1_S169: begin
        _address_addr <= 169;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S170;
      end
      retro_main_b1_S170: begin
        _address_addr <= 170;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S171;
      end
      retro_main_b1_S171: begin
        _address_addr <= 171;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S172;
      end
      retro_main_b1_S172: begin
        _address_addr <= 172;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S173;
      end
      retro_main_b1_S173: begin
        _address_addr <= 173;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S174;
      end
      retro_main_b1_S174: begin
        _address_addr <= 174;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S175;
      end
      retro_main_b1_S175: begin
        _address_addr <= 175;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S176;
      end
      retro_main_b1_S176: begin
        _address_addr <= 176;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S177;
      end
      retro_main_b1_S177: begin
        _address_addr <= 177;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S178;
      end
      retro_main_b1_S178: begin
        _address_addr <= 178;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S179;
      end
      retro_main_b1_S179: begin
        _address_addr <= 179;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S180;
      end
      retro_main_b1_S180: begin
        _address_addr <= 180;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S181;
      end
      retro_main_b1_S181: begin
        _address_addr <= 181;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S182;
      end
      retro_main_b1_S182: begin
        _address_addr <= 182;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S183;
      end
      retro_main_b1_S183: begin
        _address_addr <= 183;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S184;
      end
      retro_main_b1_S184: begin
        _address_addr <= 184;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S185;
      end
      retro_main_b1_S185: begin
        _address_addr <= 185;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S186;
      end
      retro_main_b1_S186: begin
        _address_addr <= 186;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S187;
      end
      retro_main_b1_S187: begin
        _address_addr <= 187;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S188;
      end
      retro_main_b1_S188: begin
        _address_addr <= 188;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S189;
      end
      retro_main_b1_S189: begin
        _address_addr <= 189;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S190;
      end
      retro_main_b1_S190: begin
        _address_addr <= 190;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S191;
      end
      retro_main_b1_S191: begin
        _address_addr <= 191;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S192;
      end
      retro_main_b1_S192: begin
        _address_addr <= 192;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S193;
      end
      retro_main_b1_S193: begin
        _address_addr <= 193;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S194;
      end
      retro_main_b1_S194: begin
        _address_addr <= 194;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S195;
      end
      retro_main_b1_S195: begin
        _address_addr <= 195;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S196;
      end
      retro_main_b1_S196: begin
        _address_addr <= 196;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S197;
      end
      retro_main_b1_S197: begin
        _address_addr <= 197;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S198;
      end
      retro_main_b1_S198: begin
        _address_addr <= 198;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S199;
      end
      retro_main_b1_S199: begin
        _address_addr <= 199;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S200;
      end
      retro_main_b1_S200: begin
        _address_addr <= 200;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S201;
      end
      retro_main_b1_S201: begin
        _address_addr <= 201;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S202;
      end
      retro_main_b1_S202: begin
        _address_addr <= 202;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S203;
      end
      retro_main_b1_S203: begin
        _address_addr <= 203;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S204;
      end
      retro_main_b1_S204: begin
        _address_addr <= 204;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S205;
      end
      retro_main_b1_S205: begin
        _address_addr <= 205;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S206;
      end
      retro_main_b1_S206: begin
        _address_addr <= 206;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S207;
      end
      retro_main_b1_S207: begin
        _address_addr <= 207;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S208;
      end
      retro_main_b1_S208: begin
        _address_addr <= 208;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S209;
      end
      retro_main_b1_S209: begin
        _address_addr <= 209;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S210;
      end
      retro_main_b1_S210: begin
        _address_addr <= 210;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S211;
      end
      retro_main_b1_S211: begin
        _address_addr <= 211;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S212;
      end
      retro_main_b1_S212: begin
        _address_addr <= 212;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S213;
      end
      retro_main_b1_S213: begin
        _address_addr <= 213;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S214;
      end
      retro_main_b1_S214: begin
        _address_addr <= 214;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S215;
      end
      retro_main_b1_S215: begin
        _address_addr <= 215;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S216;
      end
      retro_main_b1_S216: begin
        _address_addr <= 216;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S217;
      end
      retro_main_b1_S217: begin
        _address_addr <= 217;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S218;
      end
      retro_main_b1_S218: begin
        _address_addr <= 218;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S219;
      end
      retro_main_b1_S219: begin
        _address_addr <= 219;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S220;
      end
      retro_main_b1_S220: begin
        _address_addr <= 220;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S221;
      end
      retro_main_b1_S221: begin
        _address_addr <= 221;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S222;
      end
      retro_main_b1_S222: begin
        _address_addr <= 222;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S223;
      end
      retro_main_b1_S223: begin
        _address_addr <= 223;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S224;
      end
      retro_main_b1_S224: begin
        _address_addr <= 224;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S225;
      end
      retro_main_b1_S225: begin
        _address_addr <= 225;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S226;
      end
      retro_main_b1_S226: begin
        _address_addr <= 226;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S227;
      end
      retro_main_b1_S227: begin
        _address_addr <= 227;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S228;
      end
      retro_main_b1_S228: begin
        _address_addr <= 228;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S229;
      end
      retro_main_b1_S229: begin
        _address_addr <= 229;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S230;
      end
      retro_main_b1_S230: begin
        _address_addr <= 230;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S231;
      end
      retro_main_b1_S231: begin
        _address_addr <= 231;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S232;
      end
      retro_main_b1_S232: begin
        _address_addr <= 232;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S233;
      end
      retro_main_b1_S233: begin
        _address_addr <= 233;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S234;
      end
      retro_main_b1_S234: begin
        _address_addr <= 234;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S235;
      end
      retro_main_b1_S235: begin
        _address_addr <= 235;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S236;
      end
      retro_main_b1_S236: begin
        _address_addr <= 236;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S237;
      end
      retro_main_b1_S237: begin
        _address_addr <= 237;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S238;
      end
      retro_main_b1_S238: begin
        _address_addr <= 238;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S239;
      end
      retro_main_b1_S239: begin
        _address_addr <= 239;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S240;
      end
      retro_main_b1_S240: begin
        _address_addr <= 240;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S241;
      end
      retro_main_b1_S241: begin
        _address_addr <= 241;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S242;
      end
      retro_main_b1_S242: begin
        _address_addr <= 242;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S243;
      end
      retro_main_b1_S243: begin
        _address_addr <= 243;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S244;
      end
      retro_main_b1_S244: begin
        _address_addr <= 244;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S245;
      end
      retro_main_b1_S245: begin
        _address_addr <= 245;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S246;
      end
      retro_main_b1_S246: begin
        _address_addr <= 246;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S247;
      end
      retro_main_b1_S247: begin
        _address_addr <= 247;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S248;
      end
      retro_main_b1_S248: begin
        _address_addr <= 248;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S249;
      end
      retro_main_b1_S249: begin
        _address_addr <= 249;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S250;
      end
      retro_main_b1_S250: begin
        _address_addr <= 250;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S251;
      end
      retro_main_b1_S251: begin
        _address_addr <= 251;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S252;
      end
      retro_main_b1_S252: begin
        _address_addr <= 252;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S253;
      end
      retro_main_b1_S253: begin
        _address_addr <= 253;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S254;
      end
      retro_main_b1_S254: begin
        _address_addr <= 254;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S255;
      end
      retro_main_b1_S255: begin
        _address_addr <= 255;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S256;
      end
      retro_main_b1_S256: begin
        _address_addr <= 256;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S257;
      end
      retro_main_b1_S257: begin
        _address_addr <= 257;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S258;
      end
      retro_main_b1_S258: begin
        _address_addr <= 258;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S259;
      end
      retro_main_b1_S259: begin
        _address_addr <= 259;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S260;
      end
      retro_main_b1_S260: begin
        _address_addr <= 260;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S261;
      end
      retro_main_b1_S261: begin
        _address_addr <= 261;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S262;
      end
      retro_main_b1_S262: begin
        _address_addr <= 262;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S263;
      end
      retro_main_b1_S263: begin
        _address_addr <= 263;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S264;
      end
      retro_main_b1_S264: begin
        _address_addr <= 264;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S265;
      end
      retro_main_b1_S265: begin
        _address_addr <= 265;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S266;
      end
      retro_main_b1_S266: begin
        _address_addr <= 266;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S267;
      end
      retro_main_b1_S267: begin
        _address_addr <= 267;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S268;
      end
      retro_main_b1_S268: begin
        _address_addr <= 268;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S269;
      end
      retro_main_b1_S269: begin
        _address_addr <= 269;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S270;
      end
      retro_main_b1_S270: begin
        _address_addr <= 270;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S271;
      end
      retro_main_b1_S271: begin
        _address_addr <= 271;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S272;
      end
      retro_main_b1_S272: begin
        _address_addr <= 272;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S273;
      end
      retro_main_b1_S273: begin
        _address_addr <= 273;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S274;
      end
      retro_main_b1_S274: begin
        _address_addr <= 274;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S275;
      end
      retro_main_b1_S275: begin
        _address_addr <= 275;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S276;
      end
      retro_main_b1_S276: begin
        _address_addr <= 276;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S277;
      end
      retro_main_b1_S277: begin
        _address_addr <= 277;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S278;
      end
      retro_main_b1_S278: begin
        _address_addr <= 278;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S279;
      end
      retro_main_b1_S279: begin
        _address_addr <= 279;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S280;
      end
      retro_main_b1_S280: begin
        _address_addr <= 280;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S281;
      end
      retro_main_b1_S281: begin
        _address_addr <= 281;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S282;
      end
      retro_main_b1_S282: begin
        _address_addr <= 282;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S283;
      end
      retro_main_b1_S283: begin
        _address_addr <= 283;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S284;
      end
      retro_main_b1_S284: begin
        _address_addr <= 284;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S285;
      end
      retro_main_b1_S285: begin
        _address_addr <= 285;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S286;
      end
      retro_main_b1_S286: begin
        _address_addr <= 286;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S287;
      end
      retro_main_b1_S287: begin
        _address_addr <= 287;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S288;
      end
      retro_main_b1_S288: begin
        _address_addr <= 288;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S289;
      end
      retro_main_b1_S289: begin
        _address_addr <= 289;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S290;
      end
      retro_main_b1_S290: begin
        _address_addr <= 290;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S291;
      end
      retro_main_b1_S291: begin
        _address_addr <= 291;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S292;
      end
      retro_main_b1_S292: begin
        _address_addr <= 292;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S293;
      end
      retro_main_b1_S293: begin
        _address_addr <= 293;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S294;
      end
      retro_main_b1_S294: begin
        _address_addr <= 294;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S295;
      end
      retro_main_b1_S295: begin
        _address_addr <= 295;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S296;
      end
      retro_main_b1_S296: begin
        _address_addr <= 296;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S297;
      end
      retro_main_b1_S297: begin
        _address_addr <= 297;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S298;
      end
      retro_main_b1_S298: begin
        _address_addr <= 298;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S299;
      end
      retro_main_b1_S299: begin
        _address_addr <= 299;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S300;
      end
      retro_main_b1_S300: begin
        _address_addr <= 300;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S301;
      end
      retro_main_b1_S301: begin
        _address_addr <= 301;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S302;
      end
      retro_main_b1_S302: begin
        _address_addr <= 302;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S303;
      end
      retro_main_b1_S303: begin
        _address_addr <= 303;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S304;
      end
      retro_main_b1_S304: begin
        _address_addr <= 304;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S305;
      end
      retro_main_b1_S305: begin
        _address_addr <= 305;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S306;
      end
      retro_main_b1_S306: begin
        _address_addr <= 306;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S307;
      end
      retro_main_b1_S307: begin
        _address_addr <= 307;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S308;
      end
      retro_main_b1_S308: begin
        _address_addr <= 308;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S309;
      end
      retro_main_b1_S309: begin
        _address_addr <= 309;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S310;
      end
      retro_main_b1_S310: begin
        _address_addr <= 310;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S311;
      end
      retro_main_b1_S311: begin
        _address_addr <= 311;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S312;
      end
      retro_main_b1_S312: begin
        _address_addr <= 312;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S313;
      end
      retro_main_b1_S313: begin
        _address_addr <= 313;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S314;
      end
      retro_main_b1_S314: begin
        _address_addr <= 314;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S315;
      end
      retro_main_b1_S315: begin
        _address_addr <= 315;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S316;
      end
      retro_main_b1_S316: begin
        _address_addr <= 316;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S317;
      end
      retro_main_b1_S317: begin
        _address_addr <= 317;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S318;
      end
      retro_main_b1_S318: begin
        _address_addr <= 318;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S319;
      end
      retro_main_b1_S319: begin
        _address_addr <= 319;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S320;
      end
      retro_main_b1_S320: begin
        _address_addr <= 320;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S321;
      end
      retro_main_b1_S321: begin
        _address_addr <= 321;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S322;
      end
      retro_main_b1_S322: begin
        _address_addr <= 322;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S323;
      end
      retro_main_b1_S323: begin
        _address_addr <= 323;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S324;
      end
      retro_main_b1_S324: begin
        _address_addr <= 324;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S325;
      end
      retro_main_b1_S325: begin
        _address_addr <= 325;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S326;
      end
      retro_main_b1_S326: begin
        _address_addr <= 326;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S327;
      end
      retro_main_b1_S327: begin
        _address_addr <= 327;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S328;
      end
      retro_main_b1_S328: begin
        _address_addr <= 328;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S329;
      end
      retro_main_b1_S329: begin
        _address_addr <= 329;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S330;
      end
      retro_main_b1_S330: begin
        _address_addr <= 330;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S331;
      end
      retro_main_b1_S331: begin
        _address_addr <= 331;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S332;
      end
      retro_main_b1_S332: begin
        _address_addr <= 332;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S333;
      end
      retro_main_b1_S333: begin
        _address_addr <= 333;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S334;
      end
      retro_main_b1_S334: begin
        _address_addr <= 334;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S335;
      end
      retro_main_b1_S335: begin
        _address_addr <= 335;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S336;
      end
      retro_main_b1_S336: begin
        _address_addr <= 336;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S337;
      end
      retro_main_b1_S337: begin
        _address_addr <= 337;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S338;
      end
      retro_main_b1_S338: begin
        _address_addr <= 338;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S339;
      end
      retro_main_b1_S339: begin
        _address_addr <= 339;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S340;
      end
      retro_main_b1_S340: begin
        _address_addr <= 340;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S341;
      end
      retro_main_b1_S341: begin
        _address_addr <= 341;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S342;
      end
      retro_main_b1_S342: begin
        _address_addr <= 342;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S343;
      end
      retro_main_b1_S343: begin
        _address_addr <= 343;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S344;
      end
      retro_main_b1_S344: begin
        _address_addr <= 344;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S345;
      end
      retro_main_b1_S345: begin
        _address_addr <= 345;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S346;
      end
      retro_main_b1_S346: begin
        _address_addr <= 346;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S347;
      end
      retro_main_b1_S347: begin
        _address_addr <= 347;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S348;
      end
      retro_main_b1_S348: begin
        _address_addr <= 348;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S349;
      end
      retro_main_b1_S349: begin
        _address_addr <= 349;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S350;
      end
      retro_main_b1_S350: begin
        _address_addr <= 350;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S351;
      end
      retro_main_b1_S351: begin
        _address_addr <= 351;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S352;
      end
      retro_main_b1_S352: begin
        _address_addr <= 352;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S353;
      end
      retro_main_b1_S353: begin
        _address_addr <= 353;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S354;
      end
      retro_main_b1_S354: begin
        _address_addr <= 354;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S355;
      end
      retro_main_b1_S355: begin
        _address_addr <= 355;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S356;
      end
      retro_main_b1_S356: begin
        _address_addr <= 356;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S357;
      end
      retro_main_b1_S357: begin
        _address_addr <= 357;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S358;
      end
      retro_main_b1_S358: begin
        _address_addr <= 358;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S359;
      end
      retro_main_b1_S359: begin
        _address_addr <= 359;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S360;
      end
      retro_main_b1_S360: begin
        _address_addr <= 360;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S361;
      end
      retro_main_b1_S361: begin
        _address_addr <= 361;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S362;
      end
      retro_main_b1_S362: begin
        _address_addr <= 362;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S363;
      end
      retro_main_b1_S363: begin
        _address_addr <= 363;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S364;
      end
      retro_main_b1_S364: begin
        _address_addr <= 364;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S365;
      end
      retro_main_b1_S365: begin
        _address_addr <= 365;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S366;
      end
      retro_main_b1_S366: begin
        _address_addr <= 366;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S367;
      end
      retro_main_b1_S367: begin
        _address_addr <= 367;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S368;
      end
      retro_main_b1_S368: begin
        _address_addr <= 368;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S369;
      end
      retro_main_b1_S369: begin
        _address_addr <= 369;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S370;
      end
      retro_main_b1_S370: begin
        _address_addr <= 370;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S371;
      end
      retro_main_b1_S371: begin
        _address_addr <= 371;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S372;
      end
      retro_main_b1_S372: begin
        _address_addr <= 372;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S373;
      end
      retro_main_b1_S373: begin
        _address_addr <= 373;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S374;
      end
      retro_main_b1_S374: begin
        _address_addr <= 374;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S375;
      end
      retro_main_b1_S375: begin
        _address_addr <= 375;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S376;
      end
      retro_main_b1_S376: begin
        _address_addr <= 376;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S377;
      end
      retro_main_b1_S377: begin
        _address_addr <= 377;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S378;
      end
      retro_main_b1_S378: begin
        _address_addr <= 378;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S379;
      end
      retro_main_b1_S379: begin
        _address_addr <= 379;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S380;
      end
      retro_main_b1_S380: begin
        _address_addr <= 380;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S381;
      end
      retro_main_b1_S381: begin
        _address_addr <= 381;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S382;
      end
      retro_main_b1_S382: begin
        _address_addr <= 382;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S383;
      end
      retro_main_b1_S383: begin
        _address_addr <= 383;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S384;
      end
      retro_main_b1_S384: begin
        _address_addr <= 384;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S385;
      end
      retro_main_b1_S385: begin
        _address_addr <= 385;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S386;
      end
      retro_main_b1_S386: begin
        _address_addr <= 386;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S387;
      end
      retro_main_b1_S387: begin
        _address_addr <= 387;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S388;
      end
      retro_main_b1_S388: begin
        _address_addr <= 388;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S389;
      end
      retro_main_b1_S389: begin
        _address_addr <= 389;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S390;
      end
      retro_main_b1_S390: begin
        _address_addr <= 390;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S391;
      end
      retro_main_b1_S391: begin
        _address_addr <= 391;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S392;
      end
      retro_main_b1_S392: begin
        _address_addr <= 392;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S393;
      end
      retro_main_b1_S393: begin
        _address_addr <= 393;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S394;
      end
      retro_main_b1_S394: begin
        _address_addr <= 394;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S395;
      end
      retro_main_b1_S395: begin
        _address_addr <= 395;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S396;
      end
      retro_main_b1_S396: begin
        _address_addr <= 396;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S397;
      end
      retro_main_b1_S397: begin
        _address_addr <= 397;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S398;
      end
      retro_main_b1_S398: begin
        _address_addr <= 398;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S399;
      end
      retro_main_b1_S399: begin
        _address_addr <= 399;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S400;
      end
      retro_main_b1_S400: begin
        _address_addr <= 400;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S401;
      end
      retro_main_b1_S401: begin
        _address_addr <= 401;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S402;
      end
      retro_main_b1_S402: begin
        _address_addr <= 402;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S403;
      end
      retro_main_b1_S403: begin
        _address_addr <= 403;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S404;
      end
      retro_main_b1_S404: begin
        _address_addr <= 404;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S405;
      end
      retro_main_b1_S405: begin
        _address_addr <= 405;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S406;
      end
      retro_main_b1_S406: begin
        _address_addr <= 406;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S407;
      end
      retro_main_b1_S407: begin
        _address_addr <= 407;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S408;
      end
      retro_main_b1_S408: begin
        _address_addr <= 408;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S409;
      end
      retro_main_b1_S409: begin
        _address_addr <= 409;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S410;
      end
      retro_main_b1_S410: begin
        _address_addr <= 410;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S411;
      end
      retro_main_b1_S411: begin
        _address_addr <= 411;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S412;
      end
      retro_main_b1_S412: begin
        _address_addr <= 412;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S413;
      end
      retro_main_b1_S413: begin
        _address_addr <= 413;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S414;
      end
      retro_main_b1_S414: begin
        _address_addr <= 414;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S415;
      end
      retro_main_b1_S415: begin
        _address_addr <= 415;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S416;
      end
      retro_main_b1_S416: begin
        _address_addr <= 416;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S417;
      end
      retro_main_b1_S417: begin
        _address_addr <= 417;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S418;
      end
      retro_main_b1_S418: begin
        _address_addr <= 418;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S419;
      end
      retro_main_b1_S419: begin
        _address_addr <= 419;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S420;
      end
      retro_main_b1_S420: begin
        _address_addr <= 420;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S421;
      end
      retro_main_b1_S421: begin
        _address_addr <= 421;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S422;
      end
      retro_main_b1_S422: begin
        _address_addr <= 422;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S423;
      end
      retro_main_b1_S423: begin
        _address_addr <= 423;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S424;
      end
      retro_main_b1_S424: begin
        _address_addr <= 424;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S425;
      end
      retro_main_b1_S425: begin
        _address_addr <= 425;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S426;
      end
      retro_main_b1_S426: begin
        _address_addr <= 426;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S427;
      end
      retro_main_b1_S427: begin
        _address_addr <= 427;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S428;
      end
      retro_main_b1_S428: begin
        _address_addr <= 428;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S429;
      end
      retro_main_b1_S429: begin
        _address_addr <= 429;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S430;
      end
      retro_main_b1_S430: begin
        _address_addr <= 430;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S431;
      end
      retro_main_b1_S431: begin
        _address_addr <= 431;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S432;
      end
      retro_main_b1_S432: begin
        _address_addr <= 432;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S433;
      end
      retro_main_b1_S433: begin
        _address_addr <= 433;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S434;
      end
      retro_main_b1_S434: begin
        _address_addr <= 434;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S435;
      end
      retro_main_b1_S435: begin
        _address_addr <= 435;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S436;
      end
      retro_main_b1_S436: begin
        _address_addr <= 436;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S437;
      end
      retro_main_b1_S437: begin
        _address_addr <= 437;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S438;
      end
      retro_main_b1_S438: begin
        _address_addr <= 438;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S439;
      end
      retro_main_b1_S439: begin
        _address_addr <= 439;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S440;
      end
      retro_main_b1_S440: begin
        _address_addr <= 440;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S441;
      end
      retro_main_b1_S441: begin
        _address_addr <= 441;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S442;
      end
      retro_main_b1_S442: begin
        _address_addr <= 442;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S443;
      end
      retro_main_b1_S443: begin
        _address_addr <= 443;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S444;
      end
      retro_main_b1_S444: begin
        _address_addr <= 444;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S445;
      end
      retro_main_b1_S445: begin
        _address_addr <= 445;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S446;
      end
      retro_main_b1_S446: begin
        _address_addr <= 446;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S447;
      end
      retro_main_b1_S447: begin
        _address_addr <= 447;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S448;
      end
      retro_main_b1_S448: begin
        _address_addr <= 448;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S449;
      end
      retro_main_b1_S449: begin
        _address_addr <= 449;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S450;
      end
      retro_main_b1_S450: begin
        _address_addr <= 450;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S451;
      end
      retro_main_b1_S451: begin
        _address_addr <= 451;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S452;
      end
      retro_main_b1_S452: begin
        _address_addr <= 452;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S453;
      end
      retro_main_b1_S453: begin
        _address_addr <= 453;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S454;
      end
      retro_main_b1_S454: begin
        _address_addr <= 454;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S455;
      end
      retro_main_b1_S455: begin
        _address_addr <= 455;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S456;
      end
      retro_main_b1_S456: begin
        _address_addr <= 456;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S457;
      end
      retro_main_b1_S457: begin
        _address_addr <= 457;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S458;
      end
      retro_main_b1_S458: begin
        _address_addr <= 458;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S459;
      end
      retro_main_b1_S459: begin
        _address_addr <= 459;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S460;
      end
      retro_main_b1_S460: begin
        _address_addr <= 460;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S461;
      end
      retro_main_b1_S461: begin
        _address_addr <= 461;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S462;
      end
      retro_main_b1_S462: begin
        _address_addr <= 462;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S463;
      end
      retro_main_b1_S463: begin
        _address_addr <= 463;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S464;
      end
      retro_main_b1_S464: begin
        _address_addr <= 464;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S465;
      end
      retro_main_b1_S465: begin
        _address_addr <= 465;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S466;
      end
      retro_main_b1_S466: begin
        _address_addr <= 466;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S467;
      end
      retro_main_b1_S467: begin
        _address_addr <= 467;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S468;
      end
      retro_main_b1_S468: begin
        _address_addr <= 468;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S469;
      end
      retro_main_b1_S469: begin
        _address_addr <= 469;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S470;
      end
      retro_main_b1_S470: begin
        _address_addr <= 470;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S471;
      end
      retro_main_b1_S471: begin
        _address_addr <= 471;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S472;
      end
      retro_main_b1_S472: begin
        _address_addr <= 472;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S473;
      end
      retro_main_b1_S473: begin
        _address_addr <= 473;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S474;
      end
      retro_main_b1_S474: begin
        _address_addr <= 474;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S475;
      end
      retro_main_b1_S475: begin
        _address_addr <= 475;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S476;
      end
      retro_main_b1_S476: begin
        _address_addr <= 476;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S477;
      end
      retro_main_b1_S477: begin
        _address_addr <= 477;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S478;
      end
      retro_main_b1_S478: begin
        _address_addr <= 478;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S479;
      end
      retro_main_b1_S479: begin
        _address_addr <= 479;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S480;
      end
      retro_main_b1_S480: begin
        _address_addr <= 480;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S481;
      end
      retro_main_b1_S481: begin
        _address_addr <= 481;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S482;
      end
      retro_main_b1_S482: begin
        _address_addr <= 482;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S483;
      end
      retro_main_b1_S483: begin
        _address_addr <= 483;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S484;
      end
      retro_main_b1_S484: begin
        _address_addr <= 484;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S485;
      end
      retro_main_b1_S485: begin
        _address_addr <= 485;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S486;
      end
      retro_main_b1_S486: begin
        _address_addr <= 486;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S487;
      end
      retro_main_b1_S487: begin
        _address_addr <= 487;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S488;
      end
      retro_main_b1_S488: begin
        _address_addr <= 488;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S489;
      end
      retro_main_b1_S489: begin
        _address_addr <= 489;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S490;
      end
      retro_main_b1_S490: begin
        _address_addr <= 490;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S491;
      end
      retro_main_b1_S491: begin
        _address_addr <= 491;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S492;
      end
      retro_main_b1_S492: begin
        _address_addr <= 492;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S493;
      end
      retro_main_b1_S493: begin
        _address_addr <= 493;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S494;
      end
      retro_main_b1_S494: begin
        _address_addr <= 494;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S495;
      end
      retro_main_b1_S495: begin
        _address_addr <= 495;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S496;
      end
      retro_main_b1_S496: begin
        _address_addr <= 496;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S497;
      end
      retro_main_b1_S497: begin
        _address_addr <= 497;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S498;
      end
      retro_main_b1_S498: begin
        _address_addr <= 498;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S499;
      end
      retro_main_b1_S499: begin
        _address_addr <= 499;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S500;
      end
      retro_main_b1_S500: begin
        _address_addr <= 500;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S501;
      end
      retro_main_b1_S501: begin
        _address_addr <= 501;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S502;
      end
      retro_main_b1_S502: begin
        _address_addr <= 502;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S503;
      end
      retro_main_b1_S503: begin
        _address_addr <= 503;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S504;
      end
      retro_main_b1_S504: begin
        _address_addr <= 504;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S505;
      end
      retro_main_b1_S505: begin
        _address_addr <= 505;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S506;
      end
      retro_main_b1_S506: begin
        _address_addr <= 506;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S507;
      end
      retro_main_b1_S507: begin
        _address_addr <= 507;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S508;
      end
      retro_main_b1_S508: begin
        _address_addr <= 508;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S509;
      end
      retro_main_b1_S509: begin
        _address_addr <= 509;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S510;
      end
      retro_main_b1_S510: begin
        _address_addr <= 510;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S511;
      end
      retro_main_b1_S511: begin
        _address_addr <= 511;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S512;
      end
      retro_main_b1_S512: begin
        _address_addr <= 512;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S513;
      end
      retro_main_b1_S513: begin
        _address_addr <= 513;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S514;
      end
      retro_main_b1_S514: begin
        _address_addr <= 514;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S515;
      end
      retro_main_b1_S515: begin
        _address_addr <= 515;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S516;
      end
      retro_main_b1_S516: begin
        _address_addr <= 516;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S517;
      end
      retro_main_b1_S517: begin
        _address_addr <= 517;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S518;
      end
      retro_main_b1_S518: begin
        _address_addr <= 518;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S519;
      end
      retro_main_b1_S519: begin
        _address_addr <= 519;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S520;
      end
      retro_main_b1_S520: begin
        _address_addr <= 520;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S521;
      end
      retro_main_b1_S521: begin
        _address_addr <= 521;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S522;
      end
      retro_main_b1_S522: begin
        _address_addr <= 522;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S523;
      end
      retro_main_b1_S523: begin
        _address_addr <= 523;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S524;
      end
      retro_main_b1_S524: begin
        _address_addr <= 524;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S525;
      end
      retro_main_b1_S525: begin
        _address_addr <= 525;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S526;
      end
      retro_main_b1_S526: begin
        _address_addr <= 526;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S527;
      end
      retro_main_b1_S527: begin
        _address_addr <= 527;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S528;
      end
      retro_main_b1_S528: begin
        _address_addr <= 528;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S529;
      end
      retro_main_b1_S529: begin
        _address_addr <= 529;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S530;
      end
      retro_main_b1_S530: begin
        _address_addr <= 530;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S531;
      end
      retro_main_b1_S531: begin
        _address_addr <= 531;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S532;
      end
      retro_main_b1_S532: begin
        _address_addr <= 532;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S533;
      end
      retro_main_b1_S533: begin
        _address_addr <= 533;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S534;
      end
      retro_main_b1_S534: begin
        _address_addr <= 534;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S535;
      end
      retro_main_b1_S535: begin
        _address_addr <= 535;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S536;
      end
      retro_main_b1_S536: begin
        _address_addr <= 536;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S537;
      end
      retro_main_b1_S537: begin
        _address_addr <= 537;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S538;
      end
      retro_main_b1_S538: begin
        _address_addr <= 538;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S539;
      end
      retro_main_b1_S539: begin
        _address_addr <= 539;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S540;
      end
      retro_main_b1_S540: begin
        _address_addr <= 540;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S541;
      end
      retro_main_b1_S541: begin
        _address_addr <= 541;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S542;
      end
      retro_main_b1_S542: begin
        _address_addr <= 542;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S543;
      end
      retro_main_b1_S543: begin
        _address_addr <= 543;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S544;
      end
      retro_main_b1_S544: begin
        _address_addr <= 544;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S545;
      end
      retro_main_b1_S545: begin
        _address_addr <= 545;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S546;
      end
      retro_main_b1_S546: begin
        _address_addr <= 546;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S547;
      end
      retro_main_b1_S547: begin
        _address_addr <= 547;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S548;
      end
      retro_main_b1_S548: begin
        _address_addr <= 548;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S549;
      end
      retro_main_b1_S549: begin
        _address_addr <= 549;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S550;
      end
      retro_main_b1_S550: begin
        _address_addr <= 550;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S551;
      end
      retro_main_b1_S551: begin
        _address_addr <= 551;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S552;
      end
      retro_main_b1_S552: begin
        _address_addr <= 552;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S553;
      end
      retro_main_b1_S553: begin
        _address_addr <= 553;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S554;
      end
      retro_main_b1_S554: begin
        _address_addr <= 554;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S555;
      end
      retro_main_b1_S555: begin
        _address_addr <= 555;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S556;
      end
      retro_main_b1_S556: begin
        _address_addr <= 556;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S557;
      end
      retro_main_b1_S557: begin
        _address_addr <= 557;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S558;
      end
      retro_main_b1_S558: begin
        _address_addr <= 558;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S559;
      end
      retro_main_b1_S559: begin
        _address_addr <= 559;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S560;
      end
      retro_main_b1_S560: begin
        _address_addr <= 560;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S561;
      end
      retro_main_b1_S561: begin
        _address_addr <= 561;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S562;
      end
      retro_main_b1_S562: begin
        _address_addr <= 562;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S563;
      end
      retro_main_b1_S563: begin
        _address_addr <= 563;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S564;
      end
      retro_main_b1_S564: begin
        _address_addr <= 564;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S565;
      end
      retro_main_b1_S565: begin
        _address_addr <= 565;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S566;
      end
      retro_main_b1_S566: begin
        _address_addr <= 566;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S567;
      end
      retro_main_b1_S567: begin
        _address_addr <= 567;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S568;
      end
      retro_main_b1_S568: begin
        _address_addr <= 568;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S569;
      end
      retro_main_b1_S569: begin
        _address_addr <= 569;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S570;
      end
      retro_main_b1_S570: begin
        _address_addr <= 570;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S571;
      end
      retro_main_b1_S571: begin
        _address_addr <= 571;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S572;
      end
      retro_main_b1_S572: begin
        _address_addr <= 572;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S573;
      end
      retro_main_b1_S573: begin
        _address_addr <= 573;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S574;
      end
      retro_main_b1_S574: begin
        _address_addr <= 574;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S575;
      end
      retro_main_b1_S575: begin
        _address_addr <= 575;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S576;
      end
      retro_main_b1_S576: begin
        _address_addr <= 576;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S577;
      end
      retro_main_b1_S577: begin
        _address_addr <= 577;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S578;
      end
      retro_main_b1_S578: begin
        _address_addr <= 578;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S579;
      end
      retro_main_b1_S579: begin
        _address_addr <= 579;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S580;
      end
      retro_main_b1_S580: begin
        _address_addr <= 580;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S581;
      end
      retro_main_b1_S581: begin
        _address_addr <= 581;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S582;
      end
      retro_main_b1_S582: begin
        _address_addr <= 582;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S583;
      end
      retro_main_b1_S583: begin
        _address_addr <= 583;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S584;
      end
      retro_main_b1_S584: begin
        _address_addr <= 584;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S585;
      end
      retro_main_b1_S585: begin
        _address_addr <= 585;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S586;
      end
      retro_main_b1_S586: begin
        _address_addr <= 586;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S587;
      end
      retro_main_b1_S587: begin
        _address_addr <= 587;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S588;
      end
      retro_main_b1_S588: begin
        _address_addr <= 588;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S589;
      end
      retro_main_b1_S589: begin
        _address_addr <= 589;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S590;
      end
      retro_main_b1_S590: begin
        _address_addr <= 590;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S591;
      end
      retro_main_b1_S591: begin
        _address_addr <= 591;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S592;
      end
      retro_main_b1_S592: begin
        _address_addr <= 592;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S593;
      end
      retro_main_b1_S593: begin
        _address_addr <= 593;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S594;
      end
      retro_main_b1_S594: begin
        _address_addr <= 594;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S595;
      end
      retro_main_b1_S595: begin
        _address_addr <= 595;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S596;
      end
      retro_main_b1_S596: begin
        _address_addr <= 596;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S597;
      end
      retro_main_b1_S597: begin
        _address_addr <= 597;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S598;
      end
      retro_main_b1_S598: begin
        _address_addr <= 598;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S599;
      end
      retro_main_b1_S599: begin
        _address_addr <= 599;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S600;
      end
      retro_main_b1_S600: begin
        _address_addr <= 600;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S601;
      end
      retro_main_b1_S601: begin
        _address_addr <= 601;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S602;
      end
      retro_main_b1_S602: begin
        _address_addr <= 602;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S603;
      end
      retro_main_b1_S603: begin
        _address_addr <= 603;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S604;
      end
      retro_main_b1_S604: begin
        _address_addr <= 604;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S605;
      end
      retro_main_b1_S605: begin
        _address_addr <= 605;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S606;
      end
      retro_main_b1_S606: begin
        _address_addr <= 606;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S607;
      end
      retro_main_b1_S607: begin
        _address_addr <= 607;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S608;
      end
      retro_main_b1_S608: begin
        _address_addr <= 608;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S609;
      end
      retro_main_b1_S609: begin
        _address_addr <= 609;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S610;
      end
      retro_main_b1_S610: begin
        _address_addr <= 610;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S611;
      end
      retro_main_b1_S611: begin
        _address_addr <= 611;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S612;
      end
      retro_main_b1_S612: begin
        _address_addr <= 612;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S613;
      end
      retro_main_b1_S613: begin
        _address_addr <= 613;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S614;
      end
      retro_main_b1_S614: begin
        _address_addr <= 614;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S615;
      end
      retro_main_b1_S615: begin
        _address_addr <= 615;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S616;
      end
      retro_main_b1_S616: begin
        _address_addr <= 616;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S617;
      end
      retro_main_b1_S617: begin
        _address_addr <= 617;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S618;
      end
      retro_main_b1_S618: begin
        _address_addr <= 618;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S619;
      end
      retro_main_b1_S619: begin
        _address_addr <= 619;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S620;
      end
      retro_main_b1_S620: begin
        _address_addr <= 620;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S621;
      end
      retro_main_b1_S621: begin
        _address_addr <= 621;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S622;
      end
      retro_main_b1_S622: begin
        _address_addr <= 622;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S623;
      end
      retro_main_b1_S623: begin
        _address_addr <= 623;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S624;
      end
      retro_main_b1_S624: begin
        _address_addr <= 624;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S625;
      end
      retro_main_b1_S625: begin
        _address_addr <= 625;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S626;
      end
      retro_main_b1_S626: begin
        _address_addr <= 626;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S627;
      end
      retro_main_b1_S627: begin
        _address_addr <= 627;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S628;
      end
      retro_main_b1_S628: begin
        _address_addr <= 628;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S629;
      end
      retro_main_b1_S629: begin
        _address_addr <= 629;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S630;
      end
      retro_main_b1_S630: begin
        _address_addr <= 630;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S631;
      end
      retro_main_b1_S631: begin
        _address_addr <= 631;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S632;
      end
      retro_main_b1_S632: begin
        _address_addr <= 632;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S633;
      end
      retro_main_b1_S633: begin
        _address_addr <= 633;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S634;
      end
      retro_main_b1_S634: begin
        _address_addr <= 634;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S635;
      end
      retro_main_b1_S635: begin
        _address_addr <= 635;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S636;
      end
      retro_main_b1_S636: begin
        _address_addr <= 636;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S637;
      end
      retro_main_b1_S637: begin
        _address_addr <= 637;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S638;
      end
      retro_main_b1_S638: begin
        _address_addr <= 638;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S639;
      end
      retro_main_b1_S639: begin
        _address_addr <= 639;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S640;
      end
      retro_main_b1_S640: begin
        _address_addr <= 640;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S641;
      end
      retro_main_b1_S641: begin
        _address_addr <= 641;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S642;
      end
      retro_main_b1_S642: begin
        _address_addr <= 642;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S643;
      end
      retro_main_b1_S643: begin
        _address_addr <= 643;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S644;
      end
      retro_main_b1_S644: begin
        _address_addr <= 644;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S645;
      end
      retro_main_b1_S645: begin
        _address_addr <= 645;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S646;
      end
      retro_main_b1_S646: begin
        _address_addr <= 646;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S647;
      end
      retro_main_b1_S647: begin
        _address_addr <= 647;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S648;
      end
      retro_main_b1_S648: begin
        _address_addr <= 648;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S649;
      end
      retro_main_b1_S649: begin
        _address_addr <= 649;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S650;
      end
      retro_main_b1_S650: begin
        _address_addr <= 650;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S651;
      end
      retro_main_b1_S651: begin
        _address_addr <= 651;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S652;
      end
      retro_main_b1_S652: begin
        _address_addr <= 652;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S653;
      end
      retro_main_b1_S653: begin
        _address_addr <= 653;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S654;
      end
      retro_main_b1_S654: begin
        _address_addr <= 654;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S655;
      end
      retro_main_b1_S655: begin
        _address_addr <= 655;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S656;
      end
      retro_main_b1_S656: begin
        _address_addr <= 656;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S657;
      end
      retro_main_b1_S657: begin
        _address_addr <= 657;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S658;
      end
      retro_main_b1_S658: begin
        _address_addr <= 658;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S659;
      end
      retro_main_b1_S659: begin
        _address_addr <= 659;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S660;
      end
      retro_main_b1_S660: begin
        _address_addr <= 660;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S661;
      end
      retro_main_b1_S661: begin
        _address_addr <= 661;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S662;
      end
      retro_main_b1_S662: begin
        _address_addr <= 662;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S663;
      end
      retro_main_b1_S663: begin
        _address_addr <= 663;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S664;
      end
      retro_main_b1_S664: begin
        _address_addr <= 664;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S665;
      end
      retro_main_b1_S665: begin
        _address_addr <= 665;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S666;
      end
      retro_main_b1_S666: begin
        _address_addr <= 666;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S667;
      end
      retro_main_b1_S667: begin
        _address_addr <= 667;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S668;
      end
      retro_main_b1_S668: begin
        _address_addr <= 668;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S669;
      end
      retro_main_b1_S669: begin
        _address_addr <= 669;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S670;
      end
      retro_main_b1_S670: begin
        _address_addr <= 670;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S671;
      end
      retro_main_b1_S671: begin
        _address_addr <= 671;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S672;
      end
      retro_main_b1_S672: begin
        _address_addr <= 672;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S673;
      end
      retro_main_b1_S673: begin
        _address_addr <= 673;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S674;
      end
      retro_main_b1_S674: begin
        _address_addr <= 674;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S675;
      end
      retro_main_b1_S675: begin
        _address_addr <= 675;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S676;
      end
      retro_main_b1_S676: begin
        _address_addr <= 676;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S677;
      end
      retro_main_b1_S677: begin
        _address_addr <= 677;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S678;
      end
      retro_main_b1_S678: begin
        _address_addr <= 678;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S679;
      end
      retro_main_b1_S679: begin
        _address_addr <= 679;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S680;
      end
      retro_main_b1_S680: begin
        _address_addr <= 680;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S681;
      end
      retro_main_b1_S681: begin
        _address_addr <= 681;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S682;
      end
      retro_main_b1_S682: begin
        _address_addr <= 682;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S683;
      end
      retro_main_b1_S683: begin
        _address_addr <= 683;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S684;
      end
      retro_main_b1_S684: begin
        _address_addr <= 684;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S685;
      end
      retro_main_b1_S685: begin
        _address_addr <= 685;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S686;
      end
      retro_main_b1_S686: begin
        _address_addr <= 686;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S687;
      end
      retro_main_b1_S687: begin
        _address_addr <= 687;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S688;
      end
      retro_main_b1_S688: begin
        _address_addr <= 688;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S689;
      end
      retro_main_b1_S689: begin
        _address_addr <= 689;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S690;
      end
      retro_main_b1_S690: begin
        _address_addr <= 690;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S691;
      end
      retro_main_b1_S691: begin
        _address_addr <= 691;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S692;
      end
      retro_main_b1_S692: begin
        _address_addr <= 692;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S693;
      end
      retro_main_b1_S693: begin
        _address_addr <= 693;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S694;
      end
      retro_main_b1_S694: begin
        _address_addr <= 694;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S695;
      end
      retro_main_b1_S695: begin
        _address_addr <= 695;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S696;
      end
      retro_main_b1_S696: begin
        _address_addr <= 696;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S697;
      end
      retro_main_b1_S697: begin
        _address_addr <= 697;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S698;
      end
      retro_main_b1_S698: begin
        _address_addr <= 698;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S699;
      end
      retro_main_b1_S699: begin
        _address_addr <= 699;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S700;
      end
      retro_main_b1_S700: begin
        _address_addr <= 700;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S701;
      end
      retro_main_b1_S701: begin
        _address_addr <= 701;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S702;
      end
      retro_main_b1_S702: begin
        _address_addr <= 702;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S703;
      end
      retro_main_b1_S703: begin
        _address_addr <= 703;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S704;
      end
      retro_main_b1_S704: begin
        _address_addr <= 704;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S705;
      end
      retro_main_b1_S705: begin
        _address_addr <= 705;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S706;
      end
      retro_main_b1_S706: begin
        _address_addr <= 706;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S707;
      end
      retro_main_b1_S707: begin
        _address_addr <= 707;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S708;
      end
      retro_main_b1_S708: begin
        _address_addr <= 708;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S709;
      end
      retro_main_b1_S709: begin
        _address_addr <= 709;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S710;
      end
      retro_main_b1_S710: begin
        _address_addr <= 710;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S711;
      end
      retro_main_b1_S711: begin
        _address_addr <= 711;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S712;
      end
      retro_main_b1_S712: begin
        _address_addr <= 712;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S713;
      end
      retro_main_b1_S713: begin
        _address_addr <= 713;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S714;
      end
      retro_main_b1_S714: begin
        _address_addr <= 714;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S715;
      end
      retro_main_b1_S715: begin
        _address_addr <= 715;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S716;
      end
      retro_main_b1_S716: begin
        _address_addr <= 716;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S717;
      end
      retro_main_b1_S717: begin
        _address_addr <= 717;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S718;
      end
      retro_main_b1_S718: begin
        _address_addr <= 718;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S719;
      end
      retro_main_b1_S719: begin
        _address_addr <= 719;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S720;
      end
      retro_main_b1_S720: begin
        _address_addr <= 720;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S721;
      end
      retro_main_b1_S721: begin
        _address_addr <= 721;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S722;
      end
      retro_main_b1_S722: begin
        _address_addr <= 722;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S723;
      end
      retro_main_b1_S723: begin
        _address_addr <= 723;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S724;
      end
      retro_main_b1_S724: begin
        _address_addr <= 724;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S725;
      end
      retro_main_b1_S725: begin
        _address_addr <= 725;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S726;
      end
      retro_main_b1_S726: begin
        _address_addr <= 726;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S727;
      end
      retro_main_b1_S727: begin
        _address_addr <= 727;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S728;
      end
      retro_main_b1_S728: begin
        _address_addr <= 728;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S729;
      end
      retro_main_b1_S729: begin
        _address_addr <= 729;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S730;
      end
      retro_main_b1_S730: begin
        _address_addr <= 730;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S731;
      end
      retro_main_b1_S731: begin
        _address_addr <= 731;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S732;
      end
      retro_main_b1_S732: begin
        _address_addr <= 732;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S733;
      end
      retro_main_b1_S733: begin
        _address_addr <= 733;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S734;
      end
      retro_main_b1_S734: begin
        _address_addr <= 734;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S735;
      end
      retro_main_b1_S735: begin
        _address_addr <= 735;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S736;
      end
      retro_main_b1_S736: begin
        _address_addr <= 736;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S737;
      end
      retro_main_b1_S737: begin
        _address_addr <= 737;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S738;
      end
      retro_main_b1_S738: begin
        _address_addr <= 738;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S739;
      end
      retro_main_b1_S739: begin
        _address_addr <= 739;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S740;
      end
      retro_main_b1_S740: begin
        _address_addr <= 740;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S741;
      end
      retro_main_b1_S741: begin
        _address_addr <= 741;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S742;
      end
      retro_main_b1_S742: begin
        _address_addr <= 742;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S743;
      end
      retro_main_b1_S743: begin
        _address_addr <= 743;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S744;
      end
      retro_main_b1_S744: begin
        _address_addr <= 744;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S745;
      end
      retro_main_b1_S745: begin
        _address_addr <= 745;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S746;
      end
      retro_main_b1_S746: begin
        _address_addr <= 746;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S747;
      end
      retro_main_b1_S747: begin
        _address_addr <= 747;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S748;
      end
      retro_main_b1_S748: begin
        _address_addr <= 748;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S749;
      end
      retro_main_b1_S749: begin
        _address_addr <= 749;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S750;
      end
      retro_main_b1_S750: begin
        _address_addr <= 750;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S751;
      end
      retro_main_b1_S751: begin
        _address_addr <= 751;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S752;
      end
      retro_main_b1_S752: begin
        _address_addr <= 752;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S753;
      end
      retro_main_b1_S753: begin
        _address_addr <= 753;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S754;
      end
      retro_main_b1_S754: begin
        _address_addr <= 754;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S755;
      end
      retro_main_b1_S755: begin
        _address_addr <= 755;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S756;
      end
      retro_main_b1_S756: begin
        _address_addr <= 756;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S757;
      end
      retro_main_b1_S757: begin
        _address_addr <= 757;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S758;
      end
      retro_main_b1_S758: begin
        _address_addr <= 758;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S759;
      end
      retro_main_b1_S759: begin
        _address_addr <= 759;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S760;
      end
      retro_main_b1_S760: begin
        _address_addr <= 760;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S761;
      end
      retro_main_b1_S761: begin
        _address_addr <= 761;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S762;
      end
      retro_main_b1_S762: begin
        _address_addr <= 762;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S763;
      end
      retro_main_b1_S763: begin
        _address_addr <= 763;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S764;
      end
      retro_main_b1_S764: begin
        _address_addr <= 764;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S765;
      end
      retro_main_b1_S765: begin
        _address_addr <= 765;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S766;
      end
      retro_main_b1_S766: begin
        _address_addr <= 766;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S767;
      end
      retro_main_b1_S767: begin
        _address_addr <= 767;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S768;
      end
      retro_main_b1_S768: begin
        _address_addr <= 768;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S769;
      end
      retro_main_b1_S769: begin
        _address_addr <= 769;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S770;
      end
      retro_main_b1_S770: begin
        _address_addr <= 770;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S771;
      end
      retro_main_b1_S771: begin
        _address_addr <= 771;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S772;
      end
      retro_main_b1_S772: begin
        _address_addr <= 772;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S773;
      end
      retro_main_b1_S773: begin
        _address_addr <= 773;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S774;
      end
      retro_main_b1_S774: begin
        _address_addr <= 774;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S775;
      end
      retro_main_b1_S775: begin
        _address_addr <= 775;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S776;
      end
      retro_main_b1_S776: begin
        _address_addr <= 776;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S777;
      end
      retro_main_b1_S777: begin
        _address_addr <= 777;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S778;
      end
      retro_main_b1_S778: begin
        _address_addr <= 778;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S779;
      end
      retro_main_b1_S779: begin
        _address_addr <= 779;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S780;
      end
      retro_main_b1_S780: begin
        _address_addr <= 780;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S781;
      end
      retro_main_b1_S781: begin
        _address_addr <= 781;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S782;
      end
      retro_main_b1_S782: begin
        _address_addr <= 782;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S783;
      end
      retro_main_b1_S783: begin
        _address_addr <= 783;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S784;
      end
      retro_main_b1_S784: begin
        _address_addr <= 784;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S785;
      end
      retro_main_b1_S785: begin
        _address_addr <= 785;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S786;
      end
      retro_main_b1_S786: begin
        _address_addr <= 786;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S787;
      end
      retro_main_b1_S787: begin
        _address_addr <= 787;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S788;
      end
      retro_main_b1_S788: begin
        _address_addr <= 788;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S789;
      end
      retro_main_b1_S789: begin
        _address_addr <= 789;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S790;
      end
      retro_main_b1_S790: begin
        _address_addr <= 790;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S791;
      end
      retro_main_b1_S791: begin
        _address_addr <= 791;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S792;
      end
      retro_main_b1_S792: begin
        _address_addr <= 792;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S793;
      end
      retro_main_b1_S793: begin
        _address_addr <= 793;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S794;
      end
      retro_main_b1_S794: begin
        _address_addr <= 794;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S795;
      end
      retro_main_b1_S795: begin
        _address_addr <= 795;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S796;
      end
      retro_main_b1_S796: begin
        _address_addr <= 796;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S797;
      end
      retro_main_b1_S797: begin
        _address_addr <= 797;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S798;
      end
      retro_main_b1_S798: begin
        _address_addr <= 798;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S799;
      end
      retro_main_b1_S799: begin
        _address_addr <= 799;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S800;
      end
      retro_main_b1_S800: begin
        _address_addr <= 800;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S801;
      end
      retro_main_b1_S801: begin
        _address_addr <= 801;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S802;
      end
      retro_main_b1_S802: begin
        _address_addr <= 802;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S803;
      end
      retro_main_b1_S803: begin
        _address_addr <= 803;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S804;
      end
      retro_main_b1_S804: begin
        _address_addr <= 804;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S805;
      end
      retro_main_b1_S805: begin
        _address_addr <= 805;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S806;
      end
      retro_main_b1_S806: begin
        _address_addr <= 806;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S807;
      end
      retro_main_b1_S807: begin
        _address_addr <= 807;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S808;
      end
      retro_main_b1_S808: begin
        _address_addr <= 808;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S809;
      end
      retro_main_b1_S809: begin
        _address_addr <= 809;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S810;
      end
      retro_main_b1_S810: begin
        _address_addr <= 810;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S811;
      end
      retro_main_b1_S811: begin
        _address_addr <= 811;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S812;
      end
      retro_main_b1_S812: begin
        _address_addr <= 812;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S813;
      end
      retro_main_b1_S813: begin
        _address_addr <= 813;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S814;
      end
      retro_main_b1_S814: begin
        _address_addr <= 814;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S815;
      end
      retro_main_b1_S815: begin
        _address_addr <= 815;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S816;
      end
      retro_main_b1_S816: begin
        _address_addr <= 816;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S817;
      end
      retro_main_b1_S817: begin
        _address_addr <= 817;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S818;
      end
      retro_main_b1_S818: begin
        _address_addr <= 818;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S819;
      end
      retro_main_b1_S819: begin
        _address_addr <= 819;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S820;
      end
      retro_main_b1_S820: begin
        _address_addr <= 820;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S821;
      end
      retro_main_b1_S821: begin
        _address_addr <= 821;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S822;
      end
      retro_main_b1_S822: begin
        _address_addr <= 822;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S823;
      end
      retro_main_b1_S823: begin
        _address_addr <= 823;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S824;
      end
      retro_main_b1_S824: begin
        _address_addr <= 824;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S825;
      end
      retro_main_b1_S825: begin
        _address_addr <= 825;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S826;
      end
      retro_main_b1_S826: begin
        _address_addr <= 826;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S827;
      end
      retro_main_b1_S827: begin
        _address_addr <= 827;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S828;
      end
      retro_main_b1_S828: begin
        _address_addr <= 828;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S829;
      end
      retro_main_b1_S829: begin
        _address_addr <= 829;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S830;
      end
      retro_main_b1_S830: begin
        _address_addr <= 830;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S831;
      end
      retro_main_b1_S831: begin
        _address_addr <= 831;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S832;
      end
      retro_main_b1_S832: begin
        _address_addr <= 832;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S833;
      end
      retro_main_b1_S833: begin
        _address_addr <= 833;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S834;
      end
      retro_main_b1_S834: begin
        _address_addr <= 834;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S835;
      end
      retro_main_b1_S835: begin
        _address_addr <= 835;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S836;
      end
      retro_main_b1_S836: begin
        _address_addr <= 836;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S837;
      end
      retro_main_b1_S837: begin
        _address_addr <= 837;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S838;
      end
      retro_main_b1_S838: begin
        _address_addr <= 838;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S839;
      end
      retro_main_b1_S839: begin
        _address_addr <= 839;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S840;
      end
      retro_main_b1_S840: begin
        _address_addr <= 840;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S841;
      end
      retro_main_b1_S841: begin
        _address_addr <= 841;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S842;
      end
      retro_main_b1_S842: begin
        _address_addr <= 842;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S843;
      end
      retro_main_b1_S843: begin
        _address_addr <= 843;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S844;
      end
      retro_main_b1_S844: begin
        _address_addr <= 844;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S845;
      end
      retro_main_b1_S845: begin
        _address_addr <= 845;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S846;
      end
      retro_main_b1_S846: begin
        _address_addr <= 846;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S847;
      end
      retro_main_b1_S847: begin
        _address_addr <= 847;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S848;
      end
      retro_main_b1_S848: begin
        _address_addr <= 848;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S849;
      end
      retro_main_b1_S849: begin
        _address_addr <= 849;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S850;
      end
      retro_main_b1_S850: begin
        _address_addr <= 850;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S851;
      end
      retro_main_b1_S851: begin
        _address_addr <= 851;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S852;
      end
      retro_main_b1_S852: begin
        _address_addr <= 852;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S853;
      end
      retro_main_b1_S853: begin
        _address_addr <= 853;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S854;
      end
      retro_main_b1_S854: begin
        _address_addr <= 854;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S855;
      end
      retro_main_b1_S855: begin
        _address_addr <= 855;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S856;
      end
      retro_main_b1_S856: begin
        _address_addr <= 856;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S857;
      end
      retro_main_b1_S857: begin
        _address_addr <= 857;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S858;
      end
      retro_main_b1_S858: begin
        _address_addr <= 858;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S859;
      end
      retro_main_b1_S859: begin
        _address_addr <= 859;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S860;
      end
      retro_main_b1_S860: begin
        _address_addr <= 860;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S861;
      end
      retro_main_b1_S861: begin
        _address_addr <= 861;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S862;
      end
      retro_main_b1_S862: begin
        _address_addr <= 862;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S863;
      end
      retro_main_b1_S863: begin
        _address_addr <= 863;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S864;
      end
      retro_main_b1_S864: begin
        _address_addr <= 864;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S865;
      end
      retro_main_b1_S865: begin
        _address_addr <= 865;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S866;
      end
      retro_main_b1_S866: begin
        _address_addr <= 866;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S867;
      end
      retro_main_b1_S867: begin
        _address_addr <= 867;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S868;
      end
      retro_main_b1_S868: begin
        _address_addr <= 868;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S869;
      end
      retro_main_b1_S869: begin
        _address_addr <= 869;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S870;
      end
      retro_main_b1_S870: begin
        _address_addr <= 870;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S871;
      end
      retro_main_b1_S871: begin
        _address_addr <= 871;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S872;
      end
      retro_main_b1_S872: begin
        _address_addr <= 872;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S873;
      end
      retro_main_b1_S873: begin
        _address_addr <= 873;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S874;
      end
      retro_main_b1_S874: begin
        _address_addr <= 874;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S875;
      end
      retro_main_b1_S875: begin
        _address_addr <= 875;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S876;
      end
      retro_main_b1_S876: begin
        _address_addr <= 876;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S877;
      end
      retro_main_b1_S877: begin
        _address_addr <= 877;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S878;
      end
      retro_main_b1_S878: begin
        _address_addr <= 878;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S879;
      end
      retro_main_b1_S879: begin
        _address_addr <= 879;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S880;
      end
      retro_main_b1_S880: begin
        _address_addr <= 880;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S881;
      end
      retro_main_b1_S881: begin
        _address_addr <= 881;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S882;
      end
      retro_main_b1_S882: begin
        _address_addr <= 882;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S883;
      end
      retro_main_b1_S883: begin
        _address_addr <= 883;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S884;
      end
      retro_main_b1_S884: begin
        _address_addr <= 884;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S885;
      end
      retro_main_b1_S885: begin
        _address_addr <= 885;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S886;
      end
      retro_main_b1_S886: begin
        _address_addr <= 886;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S887;
      end
      retro_main_b1_S887: begin
        _address_addr <= 887;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S888;
      end
      retro_main_b1_S888: begin
        _address_addr <= 888;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S889;
      end
      retro_main_b1_S889: begin
        _address_addr <= 889;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S890;
      end
      retro_main_b1_S890: begin
        _address_addr <= 890;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S891;
      end
      retro_main_b1_S891: begin
        _address_addr <= 891;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S892;
      end
      retro_main_b1_S892: begin
        _address_addr <= 892;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S893;
      end
      retro_main_b1_S893: begin
        _address_addr <= 893;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S894;
      end
      retro_main_b1_S894: begin
        _address_addr <= 894;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S895;
      end
      retro_main_b1_S895: begin
        _address_addr <= 895;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S896;
      end
      retro_main_b1_S896: begin
        _address_addr <= 896;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S897;
      end
      retro_main_b1_S897: begin
        _address_addr <= 897;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S898;
      end
      retro_main_b1_S898: begin
        _address_addr <= 898;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S899;
      end
      retro_main_b1_S899: begin
        _address_addr <= 899;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S900;
      end
      retro_main_b1_S900: begin
        _address_addr <= 900;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S901;
      end
      retro_main_b1_S901: begin
        _address_addr <= 901;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S902;
      end
      retro_main_b1_S902: begin
        _address_addr <= 902;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S903;
      end
      retro_main_b1_S903: begin
        _address_addr <= 903;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S904;
      end
      retro_main_b1_S904: begin
        _address_addr <= 904;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S905;
      end
      retro_main_b1_S905: begin
        _address_addr <= 905;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S906;
      end
      retro_main_b1_S906: begin
        _address_addr <= 906;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S907;
      end
      retro_main_b1_S907: begin
        _address_addr <= 907;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S908;
      end
      retro_main_b1_S908: begin
        _address_addr <= 908;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S909;
      end
      retro_main_b1_S909: begin
        _address_addr <= 909;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S910;
      end
      retro_main_b1_S910: begin
        _address_addr <= 910;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S911;
      end
      retro_main_b1_S911: begin
        _address_addr <= 911;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S912;
      end
      retro_main_b1_S912: begin
        _address_addr <= 912;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S913;
      end
      retro_main_b1_S913: begin
        _address_addr <= 913;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S914;
      end
      retro_main_b1_S914: begin
        _address_addr <= 914;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S915;
      end
      retro_main_b1_S915: begin
        _address_addr <= 915;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S916;
      end
      retro_main_b1_S916: begin
        _address_addr <= 916;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S917;
      end
      retro_main_b1_S917: begin
        _address_addr <= 917;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S918;
      end
      retro_main_b1_S918: begin
        _address_addr <= 918;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S919;
      end
      retro_main_b1_S919: begin
        _address_addr <= 919;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S920;
      end
      retro_main_b1_S920: begin
        _address_addr <= 920;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S921;
      end
      retro_main_b1_S921: begin
        _address_addr <= 921;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S922;
      end
      retro_main_b1_S922: begin
        _address_addr <= 922;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S923;
      end
      retro_main_b1_S923: begin
        _address_addr <= 923;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S924;
      end
      retro_main_b1_S924: begin
        _address_addr <= 924;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S925;
      end
      retro_main_b1_S925: begin
        _address_addr <= 925;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S926;
      end
      retro_main_b1_S926: begin
        _address_addr <= 926;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S927;
      end
      retro_main_b1_S927: begin
        _address_addr <= 927;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S928;
      end
      retro_main_b1_S928: begin
        _address_addr <= 928;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S929;
      end
      retro_main_b1_S929: begin
        _address_addr <= 929;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S930;
      end
      retro_main_b1_S930: begin
        _address_addr <= 930;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S931;
      end
      retro_main_b1_S931: begin
        _address_addr <= 931;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S932;
      end
      retro_main_b1_S932: begin
        _address_addr <= 932;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S933;
      end
      retro_main_b1_S933: begin
        _address_addr <= 933;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S934;
      end
      retro_main_b1_S934: begin
        _address_addr <= 934;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S935;
      end
      retro_main_b1_S935: begin
        _address_addr <= 935;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S936;
      end
      retro_main_b1_S936: begin
        _address_addr <= 936;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S937;
      end
      retro_main_b1_S937: begin
        _address_addr <= 937;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S938;
      end
      retro_main_b1_S938: begin
        _address_addr <= 938;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S939;
      end
      retro_main_b1_S939: begin
        _address_addr <= 939;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S940;
      end
      retro_main_b1_S940: begin
        _address_addr <= 940;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S941;
      end
      retro_main_b1_S941: begin
        _address_addr <= 941;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S942;
      end
      retro_main_b1_S942: begin
        _address_addr <= 942;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S943;
      end
      retro_main_b1_S943: begin
        _address_addr <= 943;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S944;
      end
      retro_main_b1_S944: begin
        _address_addr <= 944;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S945;
      end
      retro_main_b1_S945: begin
        _address_addr <= 945;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S946;
      end
      retro_main_b1_S946: begin
        _address_addr <= 946;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S947;
      end
      retro_main_b1_S947: begin
        _address_addr <= 947;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S948;
      end
      retro_main_b1_S948: begin
        _address_addr <= 948;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S949;
      end
      retro_main_b1_S949: begin
        _address_addr <= 949;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S950;
      end
      retro_main_b1_S950: begin
        _address_addr <= 950;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S951;
      end
      retro_main_b1_S951: begin
        _address_addr <= 951;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S952;
      end
      retro_main_b1_S952: begin
        _address_addr <= 952;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S953;
      end
      retro_main_b1_S953: begin
        _address_addr <= 953;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S954;
      end
      retro_main_b1_S954: begin
        _address_addr <= 954;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S955;
      end
      retro_main_b1_S955: begin
        _address_addr <= 955;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S956;
      end
      retro_main_b1_S956: begin
        _address_addr <= 956;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S957;
      end
      retro_main_b1_S957: begin
        _address_addr <= 957;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S958;
      end
      retro_main_b1_S958: begin
        _address_addr <= 958;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S959;
      end
      retro_main_b1_S959: begin
        _address_addr <= 959;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S960;
      end
      retro_main_b1_S960: begin
        _address_addr <= 960;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S961;
      end
      retro_main_b1_S961: begin
        _address_addr <= 961;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S962;
      end
      retro_main_b1_S962: begin
        _address_addr <= 962;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S963;
      end
      retro_main_b1_S963: begin
        _address_addr <= 963;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S964;
      end
      retro_main_b1_S964: begin
        _address_addr <= 964;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S965;
      end
      retro_main_b1_S965: begin
        _address_addr <= 965;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S966;
      end
      retro_main_b1_S966: begin
        _address_addr <= 966;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S967;
      end
      retro_main_b1_S967: begin
        _address_addr <= 967;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S968;
      end
      retro_main_b1_S968: begin
        _address_addr <= 968;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S969;
      end
      retro_main_b1_S969: begin
        _address_addr <= 969;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S970;
      end
      retro_main_b1_S970: begin
        _address_addr <= 970;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S971;
      end
      retro_main_b1_S971: begin
        _address_addr <= 971;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S972;
      end
      retro_main_b1_S972: begin
        _address_addr <= 972;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S973;
      end
      retro_main_b1_S973: begin
        _address_addr <= 973;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S974;
      end
      retro_main_b1_S974: begin
        _address_addr <= 974;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S975;
      end
      retro_main_b1_S975: begin
        _address_addr <= 975;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S976;
      end
      retro_main_b1_S976: begin
        _address_addr <= 976;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S977;
      end
      retro_main_b1_S977: begin
        _address_addr <= 977;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S978;
      end
      retro_main_b1_S978: begin
        _address_addr <= 978;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S979;
      end
      retro_main_b1_S979: begin
        _address_addr <= 979;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S980;
      end
      retro_main_b1_S980: begin
        _address_addr <= 980;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S981;
      end
      retro_main_b1_S981: begin
        _address_addr <= 981;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S982;
      end
      retro_main_b1_S982: begin
        _address_addr <= 982;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S983;
      end
      retro_main_b1_S983: begin
        _address_addr <= 983;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S984;
      end
      retro_main_b1_S984: begin
        _address_addr <= 984;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S985;
      end
      retro_main_b1_S985: begin
        _address_addr <= 985;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S986;
      end
      retro_main_b1_S986: begin
        _address_addr <= 986;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S987;
      end
      retro_main_b1_S987: begin
        _address_addr <= 987;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S988;
      end
      retro_main_b1_S988: begin
        _address_addr <= 988;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S989;
      end
      retro_main_b1_S989: begin
        _address_addr <= 989;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S990;
      end
      retro_main_b1_S990: begin
        _address_addr <= 990;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S991;
      end
      retro_main_b1_S991: begin
        _address_addr <= 991;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S992;
      end
      retro_main_b1_S992: begin
        _address_addr <= 992;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S993;
      end
      retro_main_b1_S993: begin
        _address_addr <= 993;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S994;
      end
      retro_main_b1_S994: begin
        _address_addr <= 994;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S995;
      end
      retro_main_b1_S995: begin
        _address_addr <= 995;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S996;
      end
      retro_main_b1_S996: begin
        _address_addr <= 996;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S997;
      end
      retro_main_b1_S997: begin
        _address_addr <= 997;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S998;
      end
      retro_main_b1_S998: begin
        _address_addr <= 998;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S999;
      end
      retro_main_b1_S999: begin
        _address_addr <= 999;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S1000;
      end
      retro_main_b1_S1000: begin
        _address_addr <= 1000;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S1001;
      end
      retro_main_b1_S1001: begin
        _address_addr <= 1001;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S1002;
      end
      retro_main_b1_S1002: begin
        _address_addr <= 1002;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S1003;
      end
      retro_main_b1_S1003: begin
        _address_addr <= 1003;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S1004;
      end
      retro_main_b1_S1004: begin
        _address_addr <= 1004;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S1005;
      end
      retro_main_b1_S1005: begin
        _address_addr <= 1005;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S1006;
      end
      retro_main_b1_S1006: begin
        _address_addr <= 1006;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S1007;
      end
      retro_main_b1_S1007: begin
        _address_addr <= 1007;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S1008;
      end
      retro_main_b1_S1008: begin
        _address_addr <= 1008;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S1009;
      end
      retro_main_b1_S1009: begin
        _address_addr <= 1009;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S1010;
      end
      retro_main_b1_S1010: begin
        _address_addr <= 1010;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S1011;
      end
      retro_main_b1_S1011: begin
        _address_addr <= 1011;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S1012;
      end
      retro_main_b1_S1012: begin
        _address_addr <= 1012;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S1013;
      end
      retro_main_b1_S1013: begin
        _address_addr <= 1013;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S1014;
      end
      retro_main_b1_S1014: begin
        _address_addr <= 1014;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S1015;
      end
      retro_main_b1_S1015: begin
        _address_addr <= 1015;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S1016;
      end
      retro_main_b1_S1016: begin
        _address_addr <= 1016;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S1017;
      end
      retro_main_b1_S1017: begin
        _address_addr <= 1017;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S1018;
      end
      retro_main_b1_S1018: begin
        _address_addr <= 1018;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S1019;
      end
      retro_main_b1_S1019: begin
        _address_addr <= 1019;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S1020;
      end
      retro_main_b1_S1020: begin
        _address_addr <= 1020;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S1021;
      end
      retro_main_b1_S1021: begin
        _address_addr <= 1021;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S1022;
      end
      retro_main_b1_S1022: begin
        _address_addr <= 1022;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S1023;
      end
      retro_main_b1_S1023: begin
        _address_addr <= 1023;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S1024;
      end
      retro_main_b1_S1024: begin
        _address_req <= 0;
        retro_main_state <= retro_main_L1_while2_S0;
      end
      retro_main_L1_while2_S0: begin
        /* c886 <= (ip2 < 268435455); */
        if (c886) begin
          memory_addr <= ip2;
          memory_we <= 0;
          memory_req <= 1;
          /* c887 <= (done_flag2 != 0); */
          /* c1970 <= (c886 && c887); */
          retro_main_state <= retro_main_L1_whilebody3_S1;
        end else begin
          retro_main_valid <= 1;
          if (retro_main_accept == 1) begin
            retro_main_state <= retro_main_b1_INIT;
          end
        end
      end
      retro_main_L1_whilebody3_S1: begin
        /*wait for output of memory*/
        retro_main_state <= retro_main_L1_whilebody3_S2;
      end
      retro_main_L1_whilebody3_S2: begin
        mem_data <= memory_q;
        memory_req <= 0;
        retro_main_state <= retro_main_L1_whilebody3_S3;
      end
      retro_main_L1_whilebody3_S3: begin
        /* opcode4 <= c1970 ? mem_data : (c886 && !c887) ? opcode2 : 'bz; */
        /* c888 <= (opcode4 <= 31); */
        if (c888) begin
          /* c889 <= (opcode4 == 0); */
          /* c890 <= (opcode4 == 1); */
          /* c891 <= (opcode4 == 2); */
          /* c892 <= (opcode4 == 3); */
          /* c893 <= (opcode4 == 4); */
          /* c894 <= (opcode4 == 5); */
          /* c895 <= (opcode4 == 6); */
          /* c896 <= (opcode4 == 7); */
          /* c897 <= (opcode4 == 8); */
          /* c898 <= (opcode4 == 9); */
          /* c899 <= (opcode4 == 10); */
          /* c900 <= (opcode4 == 11); */
          /* c901 <= (opcode4 == 12); */
          /* c902 <= (opcode4 == 13); */
          /* c903 <= (opcode4 == 14); */
          /* c904 <= (opcode4 == 15); */
          /* c905 <= (opcode4 == 16); */
          /* c906 <= (opcode4 == 17); */
          /* c907 <= (opcode4 == 18); */
          /* c908 <= (opcode4 == 19); */
          /* c909 <= (opcode4 == 20); */
          /* c910 <= (opcode4 == 21); */
          /* c911 <= (opcode4 == 22); */
          /* c912 <= (opcode4 == 23); */
          /* c913 <= (opcode4 == 24); */
          /* c914 <= (opcode4 == 25); */
          /* c915 <= (opcode4 == 26); */
          /* c916 <= (opcode4 == 27); */
          /* c917 <= (opcode4 == 28); */
          /* c918 <= (opcode4 == 29); */
          /* c919 <= (opcode4 == 30); */
          /* c3337 <= (c886 && c888); */
          /* c1971 <= (c886 && c888); */
          /* c1041 <= (!c889 && c890); */
          /* c1042 <= ((!c889 && !c890) && c891); */
          /* c1043 <= (((!c889 && !c890) && !c891) && c892); */
          /* c1044 <= ((((!c889 && !c890) && !c891) && !c892) && c893); */
          /* c1045 <= (((((!c889 && !c890) && !c891) && !c892) && !c893) && c894); */
          /* c1046 <= ((((((!c889 && !c890) && !c891) && !c892) && !c893) && !c894) && c895); */
          /* c1047 <= (((((((!c889 && !c890) && !c891) && !c892) && !c893) && !c894) && !c895) && c896); */
          /* c1048 <= ((((((((!c889 && !c890) && !c891) && !c892) && !c893) && !c894) && !c895) && !c896) && c897); */
          /* c1049 <= (((((((((!c889 && !c890) && !c891) && !c892) && !c893) && !c894) && !c895) && !c896) && !c897) && c898); */
          /* c1050 <= ((((((((((!c889 && !c890) && !c891) && !c892) && !c893) && !c894) && !c895) && !c896) && !c897) && !c898) && c899); */
          /* c1051 <= (((((((((((!c889 && !c890) && !c891) && !c892) && !c893) && !c894) && !c895) && !c896) && !c897) && !c898) && !c899) && c900); */
          /* c1052 <= ((((((((((((!c889 && !c890) && !c891) && !c892) && !c893) && !c894) && !c895) && !c896) && !c897) && !c898) && !c899) && !c900) && c901); */
          /* c1053 <= (((((((((((((!c889 && !c890) && !c891) && !c892) && !c893) && !c894) && !c895) && !c896) && !c897) && !c898) && !c899) && !c900) && !c901) && c902); */
          /* c1054 <= ((((((((((((((!c889 && !c890) && !c891) && !c892) && !c893) && !c894) && !c895) && !c896) && !c897) && !c898) && !c899) && !c900) && !c901) && !c902) && c903); */
          /* c1055 <= (((((((((((((((!c889 && !c890) && !c891) && !c892) && !c893) && !c894) && !c895) && !c896) && !c897) && !c898) && !c899) && !c900) && !c901) && !c902) && !c903) && c904); */
          /* c1056 <= ((((((((((((((((!c889 && !c890) && !c891) && !c892) && !c893) && !c894) && !c895) && !c896) && !c897) && !c898) && !c899) && !c900) && !c901) && !c902) && !c903) && !c904) && c905); */
          /* c1057 <= (((((((((((((((((!c889 && !c890) && !c891) && !c892) && !c893) && !c894) && !c895) && !c896) && !c897) && !c898) && !c899) && !c900) && !c901) && !c902) && !c903) && !c904) && !c905) && c906); */
          /* c1058 <= ((((((((((((((((((!c889 && !c890) && !c891) && !c892) && !c893) && !c894) && !c895) && !c896) && !c897) && !c898) && !c899) && !c900) && !c901) && !c902) && !c903) && !c904) && !c905) && !c906) && c907); */
          /* c1059 <= (((((((((((((((((((!c889 && !c890) && !c891) && !c892) && !c893) && !c894) && !c895) && !c896) && !c897) && !c898) && !c899) && !c900) && !c901) && !c902) && !c903) && !c904) && !c905) && !c906) && !c907) && c908); */
          /* c1060 <= ((((((((((((((((((((!c889 && !c890) && !c891) && !c892) && !c893) && !c894) && !c895) && !c896) && !c897) && !c898) && !c899) && !c900) && !c901) && !c902) && !c903) && !c904) && !c905) && !c906) && !c907) && !c908) && c909); */
          /* c1061 <= (((((((((((((((((((((!c889 && !c890) && !c891) && !c892) && !c893) && !c894) && !c895) && !c896) && !c897) && !c898) && !c899) && !c900) && !c901) && !c902) && !c903) && !c904) && !c905) && !c906) && !c907) && !c908) && !c909) && c910); */
          /* c1062 <= ((((((((((((((((((((((!c889 && !c890) && !c891) && !c892) && !c893) && !c894) && !c895) && !c896) && !c897) && !c898) && !c899) && !c900) && !c901) && !c902) && !c903) && !c904) && !c905) && !c906) && !c907) && !c908) && !c909) && !c910) && c911); */
          /* c1063 <= (((((((((((((((((((((((!c889 && !c890) && !c891) && !c892) && !c893) && !c894) && !c895) && !c896) && !c897) && !c898) && !c899) && !c900) && !c901) && !c902) && !c903) && !c904) && !c905) && !c906) && !c907) && !c908) && !c909) && !c910) && !c911) && c912); */
          /* c1064 <= ((((((((((((((((((((((((!c889 && !c890) && !c891) && !c892) && !c893) && !c894) && !c895) && !c896) && !c897) && !c898) && !c899) && !c900) && !c901) && !c902) && !c903) && !c904) && !c905) && !c906) && !c907) && !c908) && !c909) && !c910) && !c911) && !c912) && c913); */
          /* c1065 <= (((((((((((((((((((((((((!c889 && !c890) && !c891) && !c892) && !c893) && !c894) && !c895) && !c896) && !c897) && !c898) && !c899) && !c900) && !c901) && !c902) && !c903) && !c904) && !c905) && !c906) && !c907) && !c908) && !c909) && !c910) && !c911) && !c912) && !c913) && c914); */
          /* c1066 <= ((((((((((((((((((((((((((!c889 && !c890) && !c891) && !c892) && !c893) && !c894) && !c895) && !c896) && !c897) && !c898) && !c899) && !c900) && !c901) && !c902) && !c903) && !c904) && !c905) && !c906) && !c907) && !c908) && !c909) && !c910) && !c911) && !c912) && !c913) && !c914) && c915); */
          /* c1067 <= (((((((((((((((((((((((((((!c889 && !c890) && !c891) && !c892) && !c893) && !c894) && !c895) && !c896) && !c897) && !c898) && !c899) && !c900) && !c901) && !c902) && !c903) && !c904) && !c905) && !c906) && !c907) && !c908) && !c909) && !c910) && !c911) && !c912) && !c913) && !c914) && !c915) && c916); */
          /* c1068 <= ((((((((((((((((((((((((((((!c889 && !c890) && !c891) && !c892) && !c893) && !c894) && !c895) && !c896) && !c897) && !c898) && !c899) && !c900) && !c901) && !c902) && !c903) && !c904) && !c905) && !c906) && !c907) && !c908) && !c909) && !c910) && !c911) && !c912) && !c913) && !c914) && !c915) && !c916) && c917); */
          /* c1069 <= (((((((((((((((((((((((((((((!c889 && !c890) && !c891) && !c892) && !c893) && !c894) && !c895) && !c896) && !c897) && !c898) && !c899) && !c900) && !c901) && !c902) && !c903) && !c904) && !c905) && !c906) && !c907) && !c908) && !c909) && !c910) && !c911) && !c912) && !c913) && !c914) && !c915) && !c916) && !c917) && c918); */
          /* c1070 <= ((((((((((((((((((((((((((((((!c889 && !c890) && !c891) && !c892) && !c893) && !c894) && !c895) && !c896) && !c897) && !c898) && !c899) && !c900) && !c901) && !c902) && !c903) && !c904) && !c905) && !c906) && !c907) && !c908) && !c909) && !c910) && !c911) && !c912) && !c913) && !c914) && !c915) && !c916) && !c917) && !c918) && c919); */
          /* c1071 <= ((((((((((((((((((((((((((((((!c889 && !c890) && !c891) && !c892) && !c893) && !c894) && !c895) && !c896) && !c897) && !c898) && !c899) && !c900) && !c901) && !c902) && !c903) && !c904) && !c905) && !c906) && !c907) && !c908) && !c909) && !c910) && !c911) && !c912) && !c913) && !c914) && !c915) && !c916) && !c917) && !c918) && !c919); */
          if (c889) begin
            /* address0_pos9 <= (c1971 && c889) ? address0_pos2 : ((c2004 || c2005) || c2006) ? address0_pos2 : c1974 ? address0_pos2 : c1975 ? address0_pos2 : c1976 ? address0_pos2 : c1977 ? address0_pos3 : c1978 ? address0_pos4 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? address0_pos2 : (((c2019 || c2017) || c2018) || c2016) ? address0_pos2 : c1981 ? address0_pos5 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? address0_pos2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? address0_pos2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? address0_pos2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? address0_pos2 : (((c2038 || c2040) || c2037) || c2039) ? address0_pos2 : (c2041 || c2042) ? address0_pos2 : c1988 ? address0_pos2 : c1989 ? address0_pos2 : c1990 ? address0_pos2 : c1991 ? address0_pos2 : c1992 ? address0_pos2 : c1993 ? address0_pos2 : c1994 ? address0_pos2 : c1995 ? address0_pos2 : c1996 ? address0_pos2 : ((c2055 || c2091) || c2090) ? address0_pos7 : c1998 ? address0_pos2 : c1999 ? address0_pos2 : c2000 ? address0_pos2 : c2001 ? address0_pos2 : (c2199 || c2198) ? address0_pos2 : (c2002 && !c927) ? address0_pos2 : c1972 ? address0_pos8 : 'bz; */
            /* address0_second9 <= (c1971 && c889) ? address0_second2 : ((c2004 || c2005) || c2006) ? address0_second2 : c1974 ? address0_second2 : c1975 ? address0_second2 : c1976 ? address0_second2 : c1977 ? address0_top2 : c1978 ? address0_second4 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? address0_second2 : (((c2019 || c2017) || c2018) || c2016) ? address0_second2 : c1981 ? address0_second5 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? address0_second2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? address0_second2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? address0_second2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? address0_second2 : (((c2038 || c2040) || c2037) || c2039) ? address0_second2 : (c2041 || c2042) ? address0_second2 : c1988 ? address0_second2 : c1989 ? address0_second2 : c1990 ? address0_second2 : c1991 ? address0_second2 : c1992 ? address0_second2 : c1993 ? address0_second2 : c1994 ? address0_second2 : c1995 ? address0_second2 : c1996 ? address0_second2 : ((c2055 || c2091) || c2090) ? address0_second7 : c1998 ? address0_second2 : c1999 ? address0_second2 : c2000 ? address0_second2 : c2001 ? address0_second2 : (c2199 || c2198) ? address0_second2 : (c2002 && !c927) ? address0_second2 : c1972 ? address0_top2 : 'bz; */
            /* address0_top9 <= (c1971 && c889) ? address0_top2 : ((c2004 || c2005) || c2006) ? address0_top2 : c1974 ? address0_top2 : c1975 ? address0_top2 : c1976 ? address0_top2 : c1977 ? stack0_top2 : c1978 ? address0_second2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? address0_top2 : (((c2019 || c2017) || c2018) || c2016) ? address0_top2 : c1981 ? address0_second2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? address0_top2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? address0_top2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? address0_top2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? address0_top2 : (((c2038 || c2040) || c2037) || c2039) ? address0_top2 : (c2041 || c2042) ? address0_top2 : c1988 ? address0_top2 : c1989 ? address0_top2 : c1990 ? address0_top2 : c1991 ? address0_top2 : c1992 ? address0_top2 : c1993 ? address0_top2 : c1994 ? address0_top2 : c1995 ? address0_top2 : c1996 ? address0_top2 : ((c2055 || c2091) || c2090) ? address0_top7 : c1998 ? address0_top2 : c1999 ? address0_top2 : c2000 ? address0_top2 : c2001 ? address0_top2 : (c2199 || c2198) ? address0_top2 : (c2002 && !c927) ? address0_top2 : c1972 ? ip2 : 'bz; */
            /* done_flag13 <= (c1971 && c889) ? done_flag2 : ((c2004 || c2005) || c2006) ? exec_result135 : c1974 ? done_flag2 : c1975 ? done_flag2 : c1976 ? done_flag2 : c1977 ? done_flag2 : c1978 ? done_flag2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? exec_result336 : (((c2019 || c2017) || c2018) || c2016) ? exec_result346 : c1981 ? done_flag2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? exec_result357 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? exec_result367 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? exec_result377 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? exec_result387 : (((c2038 || c2040) || c2037) || c2039) ? exec_result396 : (c2041 || c2042) ? exec_result404 : c1988 ? done_flag2 : c1989 ? done_flag2 : c1990 ? done_flag2 : c1991 ? done_flag2 : c1992 ? done_flag2 : c1993 ? done_flag2 : c1994 ? done_flag2 : c1995 ? done_flag2 : c1996 ? done_flag2 : ((c2055 || c2091) || c2090) ? exec_result545 : c1998 ? done_flag2 : c1999 ? done_flag2 : c2000 ? done_flag2 : c2001 ? done_flag2 : (c2199 || c2198) ? done_flag2 : (c2002 && !c927) ? done_flag2 : c1972 ? done_flag2 : 'bz; */
            /* ip16 <= (c1971 && c889) ? ip2 : ((c2004 || c2005) || c2006) ? lit0_ip4 : c1974 ? ip2 : c1975 ? ip2 : c1976 ? ip2 : c1977 ? ip2 : c1978 ? ip2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? loop0_ip5 : (((c2019 || c2017) || c2018) || c2016) ? jump0_ip5 : c1981 ? address0_top2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? jump_ge0_ip5 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? jump_le0_ip5 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? jump_ne0_ip5 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? jump_eq0_ip5 : (((c2038 || c2040) || c2037) || c2039) ? point0_ip5 : (c2041 || c2042) ? write_point0_ip4 : c1988 ? ip2 : c1989 ? ip2 : c1990 ? ip2 : c1991 ? ip2 : c1992 ? ip2 : c1993 ? ip2 : c1994 ? ip2 : c1995 ? ip2 : c1996 ? ip2 : ((c2055 || c2091) || c2090) ? zero_pop_return0_ip5 : c1998 ? ip2 : c1999 ? ip2 : c2000 ? ip2 : c2001 ? ip2 : (c2199 || c2198) ? ip_inl554 : (c2002 && !c927) ? ip2 : c1972 ? ip15 : 'bz; */
            /* jump0_ip6 <= (c1971 && c889) ? jump0_ip2 : ((c2004 || c2005) || c2006) ? jump0_ip2 : c1974 ? jump0_ip2 : c1975 ? jump0_ip2 : c1976 ? jump0_ip2 : c1977 ? jump0_ip2 : c1978 ? jump0_ip2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? jump0_ip2 : (((c2019 || c2017) || c2018) || c2016) ? jump0_ip5 : c1981 ? jump0_ip2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? jump0_ip2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? jump0_ip2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? jump0_ip2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? jump0_ip2 : (((c2038 || c2040) || c2037) || c2039) ? jump0_ip2 : (c2041 || c2042) ? jump0_ip2 : c1988 ? jump0_ip2 : c1989 ? jump0_ip2 : c1990 ? jump0_ip2 : c1991 ? jump0_ip2 : c1992 ? jump0_ip2 : c1993 ? jump0_ip2 : c1994 ? jump0_ip2 : c1995 ? jump0_ip2 : c1996 ? jump0_ip2 : ((c2055 || c2091) || c2090) ? jump0_ip2 : c1998 ? jump0_ip2 : c1999 ? jump0_ip2 : c2000 ? jump0_ip2 : c2001 ? jump0_ip2 : (c2199 || c2198) ? jump0_ip2 : (c2002 && !c927) ? jump0_ip2 : c1972 ? jump0_ip2 : 'bz; */
            /* jump0_phase8 <= (c1971 && c889) ? jump0_phase2 : ((c2004 || c2005) || c2006) ? jump0_phase2 : c1974 ? jump0_phase2 : c1975 ? jump0_phase2 : c1976 ? jump0_phase2 : c1977 ? jump0_phase2 : c1978 ? jump0_phase2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? jump0_phase2 : (((c2019 || c2017) || c2018) || c2016) ? jump0_phase7 : c1981 ? jump0_phase2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? jump0_phase2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? jump0_phase2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? jump0_phase2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? jump0_phase2 : (((c2038 || c2040) || c2037) || c2039) ? jump0_phase2 : (c2041 || c2042) ? jump0_phase2 : c1988 ? jump0_phase2 : c1989 ? jump0_phase2 : c1990 ? jump0_phase2 : c1991 ? jump0_phase2 : c1992 ? jump0_phase2 : c1993 ? jump0_phase2 : c1994 ? jump0_phase2 : c1995 ? jump0_phase2 : c1996 ? jump0_phase2 : ((c2055 || c2091) || c2090) ? jump0_phase2 : c1998 ? jump0_phase2 : c1999 ? jump0_phase2 : c2000 ? jump0_phase2 : c2001 ? jump0_phase2 : (c2199 || c2198) ? jump0_phase2 : (c2002 && !c927) ? jump0_phase2 : c1972 ? jump0_phase2 : 'bz; */
            /* jump_eq0_a5 <= (c1971 && c889) ? jump_eq0_a2 : ((c2004 || c2005) || c2006) ? jump_eq0_a2 : c1974 ? jump_eq0_a2 : c1975 ? jump_eq0_a2 : c1976 ? jump_eq0_a2 : c1977 ? jump_eq0_a2 : c1978 ? jump_eq0_a2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? jump_eq0_a2 : (((c2019 || c2017) || c2018) || c2016) ? jump_eq0_a2 : c1981 ? jump_eq0_a2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? jump_eq0_a2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? jump_eq0_a2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? jump_eq0_a2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? jump_eq0_a4 : (((c2038 || c2040) || c2037) || c2039) ? jump_eq0_a2 : (c2041 || c2042) ? jump_eq0_a2 : c1988 ? jump_eq0_a2 : c1989 ? jump_eq0_a2 : c1990 ? jump_eq0_a2 : c1991 ? jump_eq0_a2 : c1992 ? jump_eq0_a2 : c1993 ? jump_eq0_a2 : c1994 ? jump_eq0_a2 : c1995 ? jump_eq0_a2 : c1996 ? jump_eq0_a2 : ((c2055 || c2091) || c2090) ? jump_eq0_a2 : c1998 ? jump_eq0_a2 : c1999 ? jump_eq0_a2 : c2000 ? jump_eq0_a2 : c2001 ? jump_eq0_a2 : (c2199 || c2198) ? jump_eq0_a2 : (c2002 && !c927) ? jump_eq0_a2 : c1972 ? jump_eq0_a2 : 'bz; */
            /* jump_eq0_ip6 <= (c1971 && c889) ? jump_eq0_ip2 : ((c2004 || c2005) || c2006) ? jump_eq0_ip2 : c1974 ? jump_eq0_ip2 : c1975 ? jump_eq0_ip2 : c1976 ? jump_eq0_ip2 : c1977 ? jump_eq0_ip2 : c1978 ? jump_eq0_ip2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? jump_eq0_ip2 : (((c2019 || c2017) || c2018) || c2016) ? jump_eq0_ip2 : c1981 ? jump_eq0_ip2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? jump_eq0_ip2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? jump_eq0_ip2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? jump_eq0_ip2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? jump_eq0_ip5 : (((c2038 || c2040) || c2037) || c2039) ? jump_eq0_ip2 : (c2041 || c2042) ? jump_eq0_ip2 : c1988 ? jump_eq0_ip2 : c1989 ? jump_eq0_ip2 : c1990 ? jump_eq0_ip2 : c1991 ? jump_eq0_ip2 : c1992 ? jump_eq0_ip2 : c1993 ? jump_eq0_ip2 : c1994 ? jump_eq0_ip2 : c1995 ? jump_eq0_ip2 : c1996 ? jump_eq0_ip2 : ((c2055 || c2091) || c2090) ? jump_eq0_ip2 : c1998 ? jump_eq0_ip2 : c1999 ? jump_eq0_ip2 : c2000 ? jump_eq0_ip2 : c2001 ? jump_eq0_ip2 : (c2199 || c2198) ? jump_eq0_ip2 : (c2002 && !c927) ? jump_eq0_ip2 : c1972 ? jump_eq0_ip2 : 'bz; */
            /* jump_eq0_phase9 <= (c1971 && c889) ? jump_eq0_phase2 : ((c2004 || c2005) || c2006) ? jump_eq0_phase2 : c1974 ? jump_eq0_phase2 : c1975 ? jump_eq0_phase2 : c1976 ? jump_eq0_phase2 : c1977 ? jump_eq0_phase2 : c1978 ? jump_eq0_phase2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? jump_eq0_phase2 : (((c2019 || c2017) || c2018) || c2016) ? jump_eq0_phase2 : c1981 ? jump_eq0_phase2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? jump_eq0_phase2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? jump_eq0_phase2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? jump_eq0_phase2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? jump_eq0_phase8 : (((c2038 || c2040) || c2037) || c2039) ? jump_eq0_phase2 : (c2041 || c2042) ? jump_eq0_phase2 : c1988 ? jump_eq0_phase2 : c1989 ? jump_eq0_phase2 : c1990 ? jump_eq0_phase2 : c1991 ? jump_eq0_phase2 : c1992 ? jump_eq0_phase2 : c1993 ? jump_eq0_phase2 : c1994 ? jump_eq0_phase2 : c1995 ? jump_eq0_phase2 : c1996 ? jump_eq0_phase2 : ((c2055 || c2091) || c2090) ? jump_eq0_phase2 : c1998 ? jump_eq0_phase2 : c1999 ? jump_eq0_phase2 : c2000 ? jump_eq0_phase2 : c2001 ? jump_eq0_phase2 : (c2199 || c2198) ? jump_eq0_phase2 : (c2002 && !c927) ? jump_eq0_phase2 : c1972 ? jump_eq0_phase2 : 'bz; */
            /* jump_ge0_a5 <= (c1971 && c889) ? jump_ge0_a2 : ((c2004 || c2005) || c2006) ? jump_ge0_a2 : c1974 ? jump_ge0_a2 : c1975 ? jump_ge0_a2 : c1976 ? jump_ge0_a2 : c1977 ? jump_ge0_a2 : c1978 ? jump_ge0_a2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? jump_ge0_a2 : (((c2019 || c2017) || c2018) || c2016) ? jump_ge0_a2 : c1981 ? jump_ge0_a2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? jump_ge0_a4 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? jump_ge0_a2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? jump_ge0_a2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? jump_ge0_a2 : (((c2038 || c2040) || c2037) || c2039) ? jump_ge0_a2 : (c2041 || c2042) ? jump_ge0_a2 : c1988 ? jump_ge0_a2 : c1989 ? jump_ge0_a2 : c1990 ? jump_ge0_a2 : c1991 ? jump_ge0_a2 : c1992 ? jump_ge0_a2 : c1993 ? jump_ge0_a2 : c1994 ? jump_ge0_a2 : c1995 ? jump_ge0_a2 : c1996 ? jump_ge0_a2 : ((c2055 || c2091) || c2090) ? jump_ge0_a2 : c1998 ? jump_ge0_a2 : c1999 ? jump_ge0_a2 : c2000 ? jump_ge0_a2 : c2001 ? jump_ge0_a2 : (c2199 || c2198) ? jump_ge0_a2 : (c2002 && !c927) ? jump_ge0_a2 : c1972 ? jump_ge0_a2 : 'bz; */
            /* jump_ge0_ip6 <= (c1971 && c889) ? jump_ge0_ip2 : ((c2004 || c2005) || c2006) ? jump_ge0_ip2 : c1974 ? jump_ge0_ip2 : c1975 ? jump_ge0_ip2 : c1976 ? jump_ge0_ip2 : c1977 ? jump_ge0_ip2 : c1978 ? jump_ge0_ip2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? jump_ge0_ip2 : (((c2019 || c2017) || c2018) || c2016) ? jump_ge0_ip2 : c1981 ? jump_ge0_ip2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? jump_ge0_ip5 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? jump_ge0_ip2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? jump_ge0_ip2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? jump_ge0_ip2 : (((c2038 || c2040) || c2037) || c2039) ? jump_ge0_ip2 : (c2041 || c2042) ? jump_ge0_ip2 : c1988 ? jump_ge0_ip2 : c1989 ? jump_ge0_ip2 : c1990 ? jump_ge0_ip2 : c1991 ? jump_ge0_ip2 : c1992 ? jump_ge0_ip2 : c1993 ? jump_ge0_ip2 : c1994 ? jump_ge0_ip2 : c1995 ? jump_ge0_ip2 : c1996 ? jump_ge0_ip2 : ((c2055 || c2091) || c2090) ? jump_ge0_ip2 : c1998 ? jump_ge0_ip2 : c1999 ? jump_ge0_ip2 : c2000 ? jump_ge0_ip2 : c2001 ? jump_ge0_ip2 : (c2199 || c2198) ? jump_ge0_ip2 : (c2002 && !c927) ? jump_ge0_ip2 : c1972 ? jump_ge0_ip2 : 'bz; */
            /* jump_ge0_phase9 <= (c1971 && c889) ? jump_ge0_phase2 : ((c2004 || c2005) || c2006) ? jump_ge0_phase2 : c1974 ? jump_ge0_phase2 : c1975 ? jump_ge0_phase2 : c1976 ? jump_ge0_phase2 : c1977 ? jump_ge0_phase2 : c1978 ? jump_ge0_phase2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? jump_ge0_phase2 : (((c2019 || c2017) || c2018) || c2016) ? jump_ge0_phase2 : c1981 ? jump_ge0_phase2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? jump_ge0_phase8 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? jump_ge0_phase2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? jump_ge0_phase2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? jump_ge0_phase2 : (((c2038 || c2040) || c2037) || c2039) ? jump_ge0_phase2 : (c2041 || c2042) ? jump_ge0_phase2 : c1988 ? jump_ge0_phase2 : c1989 ? jump_ge0_phase2 : c1990 ? jump_ge0_phase2 : c1991 ? jump_ge0_phase2 : c1992 ? jump_ge0_phase2 : c1993 ? jump_ge0_phase2 : c1994 ? jump_ge0_phase2 : c1995 ? jump_ge0_phase2 : c1996 ? jump_ge0_phase2 : ((c2055 || c2091) || c2090) ? jump_ge0_phase2 : c1998 ? jump_ge0_phase2 : c1999 ? jump_ge0_phase2 : c2000 ? jump_ge0_phase2 : c2001 ? jump_ge0_phase2 : (c2199 || c2198) ? jump_ge0_phase2 : (c2002 && !c927) ? jump_ge0_phase2 : c1972 ? jump_ge0_phase2 : 'bz; */
            /* jump_le0_a5 <= (c1971 && c889) ? jump_le0_a2 : ((c2004 || c2005) || c2006) ? jump_le0_a2 : c1974 ? jump_le0_a2 : c1975 ? jump_le0_a2 : c1976 ? jump_le0_a2 : c1977 ? jump_le0_a2 : c1978 ? jump_le0_a2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? jump_le0_a2 : (((c2019 || c2017) || c2018) || c2016) ? jump_le0_a2 : c1981 ? jump_le0_a2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? jump_le0_a2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? jump_le0_a4 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? jump_le0_a2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? jump_le0_a2 : (((c2038 || c2040) || c2037) || c2039) ? jump_le0_a2 : (c2041 || c2042) ? jump_le0_a2 : c1988 ? jump_le0_a2 : c1989 ? jump_le0_a2 : c1990 ? jump_le0_a2 : c1991 ? jump_le0_a2 : c1992 ? jump_le0_a2 : c1993 ? jump_le0_a2 : c1994 ? jump_le0_a2 : c1995 ? jump_le0_a2 : c1996 ? jump_le0_a2 : ((c2055 || c2091) || c2090) ? jump_le0_a2 : c1998 ? jump_le0_a2 : c1999 ? jump_le0_a2 : c2000 ? jump_le0_a2 : c2001 ? jump_le0_a2 : (c2199 || c2198) ? jump_le0_a2 : (c2002 && !c927) ? jump_le0_a2 : c1972 ? jump_le0_a2 : 'bz; */
            /* jump_le0_ip6 <= (c1971 && c889) ? jump_le0_ip2 : ((c2004 || c2005) || c2006) ? jump_le0_ip2 : c1974 ? jump_le0_ip2 : c1975 ? jump_le0_ip2 : c1976 ? jump_le0_ip2 : c1977 ? jump_le0_ip2 : c1978 ? jump_le0_ip2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? jump_le0_ip2 : (((c2019 || c2017) || c2018) || c2016) ? jump_le0_ip2 : c1981 ? jump_le0_ip2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? jump_le0_ip2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? jump_le0_ip5 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? jump_le0_ip2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? jump_le0_ip2 : (((c2038 || c2040) || c2037) || c2039) ? jump_le0_ip2 : (c2041 || c2042) ? jump_le0_ip2 : c1988 ? jump_le0_ip2 : c1989 ? jump_le0_ip2 : c1990 ? jump_le0_ip2 : c1991 ? jump_le0_ip2 : c1992 ? jump_le0_ip2 : c1993 ? jump_le0_ip2 : c1994 ? jump_le0_ip2 : c1995 ? jump_le0_ip2 : c1996 ? jump_le0_ip2 : ((c2055 || c2091) || c2090) ? jump_le0_ip2 : c1998 ? jump_le0_ip2 : c1999 ? jump_le0_ip2 : c2000 ? jump_le0_ip2 : c2001 ? jump_le0_ip2 : (c2199 || c2198) ? jump_le0_ip2 : (c2002 && !c927) ? jump_le0_ip2 : c1972 ? jump_le0_ip2 : 'bz; */
            /* jump_le0_phase9 <= (c1971 && c889) ? jump_le0_phase2 : ((c2004 || c2005) || c2006) ? jump_le0_phase2 : c1974 ? jump_le0_phase2 : c1975 ? jump_le0_phase2 : c1976 ? jump_le0_phase2 : c1977 ? jump_le0_phase2 : c1978 ? jump_le0_phase2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? jump_le0_phase2 : (((c2019 || c2017) || c2018) || c2016) ? jump_le0_phase2 : c1981 ? jump_le0_phase2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? jump_le0_phase2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? jump_le0_phase8 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? jump_le0_phase2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? jump_le0_phase2 : (((c2038 || c2040) || c2037) || c2039) ? jump_le0_phase2 : (c2041 || c2042) ? jump_le0_phase2 : c1988 ? jump_le0_phase2 : c1989 ? jump_le0_phase2 : c1990 ? jump_le0_phase2 : c1991 ? jump_le0_phase2 : c1992 ? jump_le0_phase2 : c1993 ? jump_le0_phase2 : c1994 ? jump_le0_phase2 : c1995 ? jump_le0_phase2 : c1996 ? jump_le0_phase2 : ((c2055 || c2091) || c2090) ? jump_le0_phase2 : c1998 ? jump_le0_phase2 : c1999 ? jump_le0_phase2 : c2000 ? jump_le0_phase2 : c2001 ? jump_le0_phase2 : (c2199 || c2198) ? jump_le0_phase2 : (c2002 && !c927) ? jump_le0_phase2 : c1972 ? jump_le0_phase2 : 'bz; */
            /* jump_ne0_a5 <= (c1971 && c889) ? jump_ne0_a2 : ((c2004 || c2005) || c2006) ? jump_ne0_a2 : c1974 ? jump_ne0_a2 : c1975 ? jump_ne0_a2 : c1976 ? jump_ne0_a2 : c1977 ? jump_ne0_a2 : c1978 ? jump_ne0_a2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? jump_ne0_a2 : (((c2019 || c2017) || c2018) || c2016) ? jump_ne0_a2 : c1981 ? jump_ne0_a2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? jump_ne0_a2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? jump_ne0_a2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? jump_ne0_a4 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? jump_ne0_a2 : (((c2038 || c2040) || c2037) || c2039) ? jump_ne0_a2 : (c2041 || c2042) ? jump_ne0_a2 : c1988 ? jump_ne0_a2 : c1989 ? jump_ne0_a2 : c1990 ? jump_ne0_a2 : c1991 ? jump_ne0_a2 : c1992 ? jump_ne0_a2 : c1993 ? jump_ne0_a2 : c1994 ? jump_ne0_a2 : c1995 ? jump_ne0_a2 : c1996 ? jump_ne0_a2 : ((c2055 || c2091) || c2090) ? jump_ne0_a2 : c1998 ? jump_ne0_a2 : c1999 ? jump_ne0_a2 : c2000 ? jump_ne0_a2 : c2001 ? jump_ne0_a2 : (c2199 || c2198) ? jump_ne0_a2 : (c2002 && !c927) ? jump_ne0_a2 : c1972 ? jump_ne0_a2 : 'bz; */
            /* jump_ne0_ip6 <= (c1971 && c889) ? jump_ne0_ip2 : ((c2004 || c2005) || c2006) ? jump_ne0_ip2 : c1974 ? jump_ne0_ip2 : c1975 ? jump_ne0_ip2 : c1976 ? jump_ne0_ip2 : c1977 ? jump_ne0_ip2 : c1978 ? jump_ne0_ip2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? jump_ne0_ip2 : (((c2019 || c2017) || c2018) || c2016) ? jump_ne0_ip2 : c1981 ? jump_ne0_ip2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? jump_ne0_ip2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? jump_ne0_ip2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? jump_ne0_ip5 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? jump_ne0_ip2 : (((c2038 || c2040) || c2037) || c2039) ? jump_ne0_ip2 : (c2041 || c2042) ? jump_ne0_ip2 : c1988 ? jump_ne0_ip2 : c1989 ? jump_ne0_ip2 : c1990 ? jump_ne0_ip2 : c1991 ? jump_ne0_ip2 : c1992 ? jump_ne0_ip2 : c1993 ? jump_ne0_ip2 : c1994 ? jump_ne0_ip2 : c1995 ? jump_ne0_ip2 : c1996 ? jump_ne0_ip2 : ((c2055 || c2091) || c2090) ? jump_ne0_ip2 : c1998 ? jump_ne0_ip2 : c1999 ? jump_ne0_ip2 : c2000 ? jump_ne0_ip2 : c2001 ? jump_ne0_ip2 : (c2199 || c2198) ? jump_ne0_ip2 : (c2002 && !c927) ? jump_ne0_ip2 : c1972 ? jump_ne0_ip2 : 'bz; */
            /* jump_ne0_phase9 <= (c1971 && c889) ? jump_ne0_phase2 : ((c2004 || c2005) || c2006) ? jump_ne0_phase2 : c1974 ? jump_ne0_phase2 : c1975 ? jump_ne0_phase2 : c1976 ? jump_ne0_phase2 : c1977 ? jump_ne0_phase2 : c1978 ? jump_ne0_phase2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? jump_ne0_phase2 : (((c2019 || c2017) || c2018) || c2016) ? jump_ne0_phase2 : c1981 ? jump_ne0_phase2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? jump_ne0_phase2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? jump_ne0_phase2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? jump_ne0_phase8 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? jump_ne0_phase2 : (((c2038 || c2040) || c2037) || c2039) ? jump_ne0_phase2 : (c2041 || c2042) ? jump_ne0_phase2 : c1988 ? jump_ne0_phase2 : c1989 ? jump_ne0_phase2 : c1990 ? jump_ne0_phase2 : c1991 ? jump_ne0_phase2 : c1992 ? jump_ne0_phase2 : c1993 ? jump_ne0_phase2 : c1994 ? jump_ne0_phase2 : c1995 ? jump_ne0_phase2 : c1996 ? jump_ne0_phase2 : ((c2055 || c2091) || c2090) ? jump_ne0_phase2 : c1998 ? jump_ne0_phase2 : c1999 ? jump_ne0_phase2 : c2000 ? jump_ne0_phase2 : c2001 ? jump_ne0_phase2 : (c2199 || c2198) ? jump_ne0_phase2 : (c2002 && !c927) ? jump_ne0_phase2 : c1972 ? jump_ne0_phase2 : 'bz; */
            /* lit0_ip5 <= (c1971 && c889) ? lit0_ip2 : ((c2004 || c2005) || c2006) ? lit0_ip4 : c1974 ? lit0_ip2 : c1975 ? lit0_ip2 : c1976 ? lit0_ip2 : c1977 ? lit0_ip2 : c1978 ? lit0_ip2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? lit0_ip2 : (((c2019 || c2017) || c2018) || c2016) ? lit0_ip2 : c1981 ? lit0_ip2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? lit0_ip2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? lit0_ip2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? lit0_ip2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? lit0_ip2 : (((c2038 || c2040) || c2037) || c2039) ? lit0_ip2 : (c2041 || c2042) ? lit0_ip2 : c1988 ? lit0_ip2 : c1989 ? lit0_ip2 : c1990 ? lit0_ip2 : c1991 ? lit0_ip2 : c1992 ? lit0_ip2 : c1993 ? lit0_ip2 : c1994 ? lit0_ip2 : c1995 ? lit0_ip2 : c1996 ? lit0_ip2 : ((c2055 || c2091) || c2090) ? lit0_ip2 : c1998 ? lit0_ip2 : c1999 ? lit0_ip2 : c2000 ? lit0_ip2 : c2001 ? lit0_ip2 : (c2199 || c2198) ? lit0_ip2 : (c2002 && !c927) ? lit0_ip2 : c1972 ? lit0_ip2 : 'bz; */
            /* lit0_phase7 <= (c1971 && c889) ? lit0_phase2 : ((c2004 || c2005) || c2006) ? lit0_phase6 : c1974 ? lit0_phase2 : c1975 ? lit0_phase2 : c1976 ? lit0_phase2 : c1977 ? lit0_phase2 : c1978 ? lit0_phase2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? lit0_phase2 : (((c2019 || c2017) || c2018) || c2016) ? lit0_phase2 : c1981 ? lit0_phase2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? lit0_phase2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? lit0_phase2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? lit0_phase2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? lit0_phase2 : (((c2038 || c2040) || c2037) || c2039) ? lit0_phase2 : (c2041 || c2042) ? lit0_phase2 : c1988 ? lit0_phase2 : c1989 ? lit0_phase2 : c1990 ? lit0_phase2 : c1991 ? lit0_phase2 : c1992 ? lit0_phase2 : c1993 ? lit0_phase2 : c1994 ? lit0_phase2 : c1995 ? lit0_phase2 : c1996 ? lit0_phase2 : ((c2055 || c2091) || c2090) ? lit0_phase2 : c1998 ? lit0_phase2 : c1999 ? lit0_phase2 : c2000 ? lit0_phase2 : c2001 ? lit0_phase2 : (c2199 || c2198) ? lit0_phase2 : (c2002 && !c927) ? lit0_phase2 : c1972 ? lit0_phase2 : 'bz; */
            /* loop0_ip6 <= (c1971 && c889) ? loop0_ip2 : ((c2004 || c2005) || c2006) ? loop0_ip2 : c1974 ? loop0_ip2 : c1975 ? loop0_ip2 : c1976 ? loop0_ip2 : c1977 ? loop0_ip2 : c1978 ? loop0_ip2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? loop0_ip5 : (((c2019 || c2017) || c2018) || c2016) ? loop0_ip2 : c1981 ? loop0_ip2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? loop0_ip2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? loop0_ip2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? loop0_ip2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? loop0_ip2 : (((c2038 || c2040) || c2037) || c2039) ? loop0_ip2 : (c2041 || c2042) ? loop0_ip2 : c1988 ? loop0_ip2 : c1989 ? loop0_ip2 : c1990 ? loop0_ip2 : c1991 ? loop0_ip2 : c1992 ? loop0_ip2 : c1993 ? loop0_ip2 : c1994 ? loop0_ip2 : c1995 ? loop0_ip2 : c1996 ? loop0_ip2 : ((c2055 || c2091) || c2090) ? loop0_ip2 : c1998 ? loop0_ip2 : c1999 ? loop0_ip2 : c2000 ? loop0_ip2 : c2001 ? loop0_ip2 : (c2199 || c2198) ? loop0_ip2 : (c2002 && !c927) ? loop0_ip2 : c1972 ? loop0_ip2 : 'bz; */
            /* loop0_phase9 <= (c1971 && c889) ? loop0_phase2 : ((c2004 || c2005) || c2006) ? loop0_phase2 : c1974 ? loop0_phase2 : c1975 ? loop0_phase2 : c1976 ? loop0_phase2 : c1977 ? loop0_phase2 : c1978 ? loop0_phase2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? loop0_phase8 : (((c2019 || c2017) || c2018) || c2016) ? loop0_phase2 : c1981 ? loop0_phase2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? loop0_phase2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? loop0_phase2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? loop0_phase2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? loop0_phase2 : (((c2038 || c2040) || c2037) || c2039) ? loop0_phase2 : (c2041 || c2042) ? loop0_phase2 : c1988 ? loop0_phase2 : c1989 ? loop0_phase2 : c1990 ? loop0_phase2 : c1991 ? loop0_phase2 : c1992 ? loop0_phase2 : c1993 ? loop0_phase2 : c1994 ? loop0_phase2 : c1995 ? loop0_phase2 : c1996 ? loop0_phase2 : ((c2055 || c2091) || c2090) ? loop0_phase2 : c1998 ? loop0_phase2 : c1999 ? loop0_phase2 : c2000 ? loop0_phase2 : c2001 ? loop0_phase2 : (c2199 || c2198) ? loop0_phase2 : (c2002 && !c927) ? loop0_phase2 : c1972 ? loop0_phase2 : 'bz; */
            /* point0_ip6 <= (c1971 && c889) ? point0_ip2 : ((c2004 || c2005) || c2006) ? point0_ip2 : c1974 ? point0_ip2 : c1975 ? point0_ip2 : c1976 ? point0_ip2 : c1977 ? point0_ip2 : c1978 ? point0_ip2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? point0_ip2 : (((c2019 || c2017) || c2018) || c2016) ? point0_ip2 : c1981 ? point0_ip2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? point0_ip2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? point0_ip2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? point0_ip2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? point0_ip2 : (((c2038 || c2040) || c2037) || c2039) ? point0_ip5 : (c2041 || c2042) ? point0_ip2 : c1988 ? point0_ip2 : c1989 ? point0_ip2 : c1990 ? point0_ip2 : c1991 ? point0_ip2 : c1992 ? point0_ip2 : c1993 ? point0_ip2 : c1994 ? point0_ip2 : c1995 ? point0_ip2 : c1996 ? point0_ip2 : ((c2055 || c2091) || c2090) ? point0_ip2 : c1998 ? point0_ip2 : c1999 ? point0_ip2 : c2000 ? point0_ip2 : c2001 ? point0_ip2 : (c2199 || c2198) ? point0_ip2 : (c2002 && !c927) ? point0_ip2 : c1972 ? point0_ip2 : 'bz; */
            /* point0_ip_saved5 <= (c1971 && c889) ? point0_ip_saved2 : ((c2004 || c2005) || c2006) ? point0_ip_saved2 : c1974 ? point0_ip_saved2 : c1975 ? point0_ip_saved2 : c1976 ? point0_ip_saved2 : c1977 ? point0_ip_saved2 : c1978 ? point0_ip_saved2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? point0_ip_saved2 : (((c2019 || c2017) || c2018) || c2016) ? point0_ip_saved2 : c1981 ? point0_ip_saved2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? point0_ip_saved2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? point0_ip_saved2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? point0_ip_saved2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? point0_ip_saved2 : (((c2038 || c2040) || c2037) || c2039) ? point0_ip_saved4 : (c2041 || c2042) ? point0_ip_saved2 : c1988 ? point0_ip_saved2 : c1989 ? point0_ip_saved2 : c1990 ? point0_ip_saved2 : c1991 ? point0_ip_saved2 : c1992 ? point0_ip_saved2 : c1993 ? point0_ip_saved2 : c1994 ? point0_ip_saved2 : c1995 ? point0_ip_saved2 : c1996 ? point0_ip_saved2 : ((c2055 || c2091) || c2090) ? point0_ip_saved2 : c1998 ? point0_ip_saved2 : c1999 ? point0_ip_saved2 : c2000 ? point0_ip_saved2 : c2001 ? point0_ip_saved2 : (c2199 || c2198) ? point0_ip_saved2 : (c2002 && !c927) ? point0_ip_saved2 : c1972 ? point0_ip_saved2 : 'bz; */
            /* point0_phase8 <= (c1971 && c889) ? point0_phase2 : ((c2004 || c2005) || c2006) ? point0_phase2 : c1974 ? point0_phase2 : c1975 ? point0_phase2 : c1976 ? point0_phase2 : c1977 ? point0_phase2 : c1978 ? point0_phase2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? point0_phase2 : (((c2019 || c2017) || c2018) || c2016) ? point0_phase2 : c1981 ? point0_phase2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? point0_phase2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? point0_phase2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? point0_phase2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? point0_phase2 : (((c2038 || c2040) || c2037) || c2039) ? point0_phase7 : (c2041 || c2042) ? point0_phase2 : c1988 ? point0_phase2 : c1989 ? point0_phase2 : c1990 ? point0_phase2 : c1991 ? point0_phase2 : c1992 ? point0_phase2 : c1993 ? point0_phase2 : c1994 ? point0_phase2 : c1995 ? point0_phase2 : c1996 ? point0_phase2 : ((c2055 || c2091) || c2090) ? point0_phase2 : c1998 ? point0_phase2 : c1999 ? point0_phase2 : c2000 ? point0_phase2 : c2001 ? point0_phase2 : (c2199 || c2198) ? point0_phase2 : (c2002 && !c927) ? point0_phase2 : c1972 ? point0_phase2 : 'bz; */
            /* stack0_pos43 <= (c1971 && c889) ? stack0_pos2 : ((c2004 || c2005) || c2006) ? stack0_pos4 : c1974 ? stack0_pos5 : c1975 ? stack0_pos6 : c1976 ? stack0_pos2 : c1977 ? stack0_pos7 : c1978 ? stack0_pos8 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? stack0_pos10 : (((c2019 || c2017) || c2018) || c2016) ? stack0_pos2 : c1981 ? stack0_pos2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? stack0_pos13 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? stack0_pos16 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? stack0_pos19 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? stack0_pos22 : (((c2038 || c2040) || c2037) || c2039) ? stack0_pos2 : (c2041 || c2042) ? stack0_pos25 : c1988 ? stack0_pos26 : c1989 ? stack0_pos27 : c1990 ? stack0_pos28 : c1991 ? stack0_pos2 : c1992 ? stack0_pos29 : c1993 ? stack0_pos30 : c1994 ? stack0_pos31 : c1995 ? stack0_pos32 : c1996 ? stack0_pos33 : ((c2055 || c2091) || c2090) ? stack0_pos35 : c1998 ? stack0_pos2 : c1999 ? stack0_pos2 : c2000 ? stack0_pos2 : c2001 ? stack0_pos37 : (c2199 || c2198) ? stack0_pos42 : (c2002 && !c927) ? stack0_pos2 : c1972 ? stack0_pos2 : 'bz; */
            /* stack0_second45 <= (c1971 && c889) ? stack0_second2 : ((c2004 || c2005) || c2006) ? stack0_second4 : c1974 ? stack0_top2 : c1975 ? stack0_second6 : c1976 ? stack0_top2 : c1977 ? stack0_second8 : c1978 ? stack0_top2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? stack0_second11 : (((c2019 || c2017) || c2018) || c2016) ? stack0_second2 : c1981 ? stack0_second2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? stack0_second14 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? stack0_second17 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? stack0_second20 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? stack0_second23 : (((c2038 || c2040) || c2037) || c2039) ? stack0_second2 : (c2041 || c2042) ? stack0_second26 : c1988 ? stack0_second27 : c1989 ? stack0_second28 : c1990 ? stack0_second29 : c1991 ? stack0_second30 : c1992 ? stack0_second31 : c1993 ? stack0_second32 : c1994 ? stack0_second33 : c1995 ? stack0_second34 : c1996 ? stack0_second35 : ((c2055 || c2091) || c2090) ? stack0_second37 : c1998 ? stack0_second2 : c1999 ? stack0_second2 : c2000 ? stack0_second2 : c2001 ? stack0_second39 : (c2199 || c2198) ? stack0_second44 : (c2002 && !c927) ? stack0_second2 : c1972 ? stack0_second2 : 'bz; */
            /* stack0_top59 <= (c1971 && c889) ? stack0_top2 : ((c2004 || c2005) || c2006) ? stack0_top4 : c1974 ? stack0_top2 : c1975 ? stack0_second2 : c1976 ? stack0_second2 : c1977 ? stack0_second2 : c1978 ? address0_top2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? stack0_top12 : (((c2019 || c2017) || c2018) || c2016) ? stack0_top2 : c1981 ? stack0_top2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? stack0_top15 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? stack0_top18 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? stack0_top21 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? stack0_top24 : (((c2038 || c2040) || c2037) || c2039) ? stack0_top26 : (c2041 || c2042) ? stack0_second2 : c1988 ? stack0_top31 : c1989 ? stack0_top33 : c1990 ? stack0_top35 : c1991 ? stack0_top36 : c1992 ? stack0_top38 : c1993 ? stack0_top40 : c1994 ? stack0_top42 : c1995 ? stack0_top44 : c1996 ? stack0_top46 : ((c2055 || c2091) || c2090) ? stack0_top48 : c1998 ? stack0_top49 : c1999 ? stack0_top50 : c2000 ? stack0_top51 : c2001 ? stack0_second38 : (c2199 || c2198) ? stack0_top58 : (c2002 && !c927) ? stack0_top2 : c1972 ? stack0_top2 : 'bz; */
            t11 <= (c1971 && c889) ? t11 : ((c2004 || c2005) || c2006) ? t11 : c1974 ? t11 : c1975 ? t11 : c1976 ? t11 : c1977 ? t11 : c1978 ? t11 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? t11 : (((c2019 || c2017) || c2018) || c2016) ? t11 : c1981 ? t11 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? t11 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? t11 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? t11 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? t11 : (((c2038 || c2040) || c2037) || c2039) ? t11 : (c2041 || c2042) ? t11 : c1988 ? stack0_top2 : c1989 ? stack0_top2 : c1990 ? stack0_top2 : c1991 ? t11 : c1992 ? stack0_top2 : c1993 ? stack0_top2 : c1994 ? stack0_top2 : c1995 ? stack0_top2 : c1996 ? stack0_top2 : ((c2055 || c2091) || c2090) ? t11 : c1998 ? t11 : c1999 ? t11 : c2000 ? stack0_top2 : c2001 ? t11 : (c2199 || c2198) ? t11 : (c2002 && !c927) ? t11 : c1972 ? t11 : 'bz;
            /* wr_flag4 <= (c1971 && c889) ? wr_flag2 : ((c2004 || c2005) || c2006) ? wr_flag2 : c1974 ? wr_flag2 : c1975 ? wr_flag2 : c1976 ? wr_flag2 : c1977 ? wr_flag2 : c1978 ? wr_flag2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? wr_flag2 : (((c2019 || c2017) || c2018) || c2016) ? wr_flag2 : c1981 ? wr_flag2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? wr_flag2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? wr_flag2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? wr_flag2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? wr_flag2 : (((c2038 || c2040) || c2037) || c2039) ? wr_flag2 : (c2041 || c2042) ? t2829 : c1988 ? wr_flag2 : c1989 ? wr_flag2 : c1990 ? wr_flag2 : c1991 ? wr_flag2 : c1992 ? wr_flag2 : c1993 ? wr_flag2 : c1994 ? wr_flag2 : c1995 ? wr_flag2 : c1996 ? wr_flag2 : ((c2055 || c2091) || c2090) ? wr_flag2 : c1998 ? wr_flag2 : c1999 ? wr_flag2 : c2000 ? wr_flag2 : c2001 ? wr_flag2 : (c2199 || c2198) ? wr_flag2 : (c2002 && !c927) ? wr_flag2 : c1972 ? wr_flag2 : 'bz; */
            /* wr_mem_addr4 <= (c1971 && c889) ? wr_mem_addr2 : ((c2004 || c2005) || c2006) ? wr_mem_addr2 : c1974 ? wr_mem_addr2 : c1975 ? wr_mem_addr2 : c1976 ? wr_mem_addr2 : c1977 ? wr_mem_addr2 : c1978 ? wr_mem_addr2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? wr_mem_addr2 : (((c2019 || c2017) || c2018) || c2016) ? wr_mem_addr2 : c1981 ? wr_mem_addr2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? wr_mem_addr2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? wr_mem_addr2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? wr_mem_addr2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? wr_mem_addr2 : (((c2038 || c2040) || c2037) || c2039) ? wr_mem_addr2 : (c2041 || c2042) ? t2830 : c1988 ? wr_mem_addr2 : c1989 ? wr_mem_addr2 : c1990 ? wr_mem_addr2 : c1991 ? wr_mem_addr2 : c1992 ? wr_mem_addr2 : c1993 ? wr_mem_addr2 : c1994 ? wr_mem_addr2 : c1995 ? wr_mem_addr2 : c1996 ? wr_mem_addr2 : ((c2055 || c2091) || c2090) ? wr_mem_addr2 : c1998 ? wr_mem_addr2 : c1999 ? wr_mem_addr2 : c2000 ? wr_mem_addr2 : c2001 ? wr_mem_addr2 : (c2199 || c2198) ? wr_mem_addr2 : (c2002 && !c927) ? wr_mem_addr2 : c1972 ? wr_mem_addr2 : 'bz; */
            /* wr_mem_data4 <= (c1971 && c889) ? wr_mem_data2 : ((c2004 || c2005) || c2006) ? wr_mem_data2 : c1974 ? wr_mem_data2 : c1975 ? wr_mem_data2 : c1976 ? wr_mem_data2 : c1977 ? wr_mem_data2 : c1978 ? wr_mem_data2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? wr_mem_data2 : (((c2019 || c2017) || c2018) || c2016) ? wr_mem_data2 : c1981 ? wr_mem_data2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? wr_mem_data2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? wr_mem_data2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? wr_mem_data2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? wr_mem_data2 : (((c2038 || c2040) || c2037) || c2039) ? wr_mem_data2 : (c2041 || c2042) ? t2831 : c1988 ? wr_mem_data2 : c1989 ? wr_mem_data2 : c1990 ? wr_mem_data2 : c1991 ? wr_mem_data2 : c1992 ? wr_mem_data2 : c1993 ? wr_mem_data2 : c1994 ? wr_mem_data2 : c1995 ? wr_mem_data2 : c1996 ? wr_mem_data2 : ((c2055 || c2091) || c2090) ? wr_mem_data2 : c1998 ? wr_mem_data2 : c1999 ? wr_mem_data2 : c2000 ? wr_mem_data2 : c2001 ? wr_mem_data2 : (c2199 || c2198) ? wr_mem_data2 : (c2002 && !c927) ? wr_mem_data2 : c1972 ? wr_mem_data2 : 'bz; */
            /* write_point0_addr5 <= (c1971 && c889) ? write_point0_addr2 : ((c2004 || c2005) || c2006) ? write_point0_addr2 : c1974 ? write_point0_addr2 : c1975 ? write_point0_addr2 : c1976 ? write_point0_addr2 : c1977 ? write_point0_addr2 : c1978 ? write_point0_addr2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? write_point0_addr2 : (((c2019 || c2017) || c2018) || c2016) ? write_point0_addr2 : c1981 ? write_point0_addr2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? write_point0_addr2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? write_point0_addr2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? write_point0_addr2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? write_point0_addr2 : (((c2038 || c2040) || c2037) || c2039) ? write_point0_addr2 : (c2041 || c2042) ? write_point0_addr4 : c1988 ? write_point0_addr2 : c1989 ? write_point0_addr2 : c1990 ? write_point0_addr2 : c1991 ? write_point0_addr2 : c1992 ? write_point0_addr2 : c1993 ? write_point0_addr2 : c1994 ? write_point0_addr2 : c1995 ? write_point0_addr2 : c1996 ? write_point0_addr2 : ((c2055 || c2091) || c2090) ? write_point0_addr2 : c1998 ? write_point0_addr2 : c1999 ? write_point0_addr2 : c2000 ? write_point0_addr2 : c2001 ? write_point0_addr2 : (c2199 || c2198) ? write_point0_addr2 : (c2002 && !c927) ? write_point0_addr2 : c1972 ? write_point0_addr2 : 'bz; */
            /* write_point0_data5 <= (c1971 && c889) ? write_point0_data2 : ((c2004 || c2005) || c2006) ? write_point0_data2 : c1974 ? write_point0_data2 : c1975 ? write_point0_data2 : c1976 ? write_point0_data2 : c1977 ? write_point0_data2 : c1978 ? write_point0_data2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? write_point0_data2 : (((c2019 || c2017) || c2018) || c2016) ? write_point0_data2 : c1981 ? write_point0_data2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? write_point0_data2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? write_point0_data2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? write_point0_data2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? write_point0_data2 : (((c2038 || c2040) || c2037) || c2039) ? write_point0_data2 : (c2041 || c2042) ? write_point0_data4 : c1988 ? write_point0_data2 : c1989 ? write_point0_data2 : c1990 ? write_point0_data2 : c1991 ? write_point0_data2 : c1992 ? write_point0_data2 : c1993 ? write_point0_data2 : c1994 ? write_point0_data2 : c1995 ? write_point0_data2 : c1996 ? write_point0_data2 : ((c2055 || c2091) || c2090) ? write_point0_data2 : c1998 ? write_point0_data2 : c1999 ? write_point0_data2 : c2000 ? write_point0_data2 : c2001 ? write_point0_data2 : (c2199 || c2198) ? write_point0_data2 : (c2002 && !c927) ? write_point0_data2 : c1972 ? write_point0_data2 : 'bz; */
            /* write_point0_ip5 <= (c1971 && c889) ? write_point0_ip2 : ((c2004 || c2005) || c2006) ? write_point0_ip2 : c1974 ? write_point0_ip2 : c1975 ? write_point0_ip2 : c1976 ? write_point0_ip2 : c1977 ? write_point0_ip2 : c1978 ? write_point0_ip2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? write_point0_ip2 : (((c2019 || c2017) || c2018) || c2016) ? write_point0_ip2 : c1981 ? write_point0_ip2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? write_point0_ip2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? write_point0_ip2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? write_point0_ip2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? write_point0_ip2 : (((c2038 || c2040) || c2037) || c2039) ? write_point0_ip2 : (c2041 || c2042) ? write_point0_ip4 : c1988 ? write_point0_ip2 : c1989 ? write_point0_ip2 : c1990 ? write_point0_ip2 : c1991 ? write_point0_ip2 : c1992 ? write_point0_ip2 : c1993 ? write_point0_ip2 : c1994 ? write_point0_ip2 : c1995 ? write_point0_ip2 : c1996 ? write_point0_ip2 : ((c2055 || c2091) || c2090) ? write_point0_ip2 : c1998 ? write_point0_ip2 : c1999 ? write_point0_ip2 : c2000 ? write_point0_ip2 : c2001 ? write_point0_ip2 : (c2199 || c2198) ? write_point0_ip2 : (c2002 && !c927) ? write_point0_ip2 : c1972 ? write_point0_ip2 : 'bz; */
            /* write_point0_phase6 <= (c1971 && c889) ? write_point0_phase2 : ((c2004 || c2005) || c2006) ? write_point0_phase2 : c1974 ? write_point0_phase2 : c1975 ? write_point0_phase2 : c1976 ? write_point0_phase2 : c1977 ? write_point0_phase2 : c1978 ? write_point0_phase2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? write_point0_phase2 : (((c2019 || c2017) || c2018) || c2016) ? write_point0_phase2 : c1981 ? write_point0_phase2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? write_point0_phase2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? write_point0_phase2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? write_point0_phase2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? write_point0_phase2 : (((c2038 || c2040) || c2037) || c2039) ? write_point0_phase2 : (c2041 || c2042) ? write_point0_phase5 : c1988 ? write_point0_phase2 : c1989 ? write_point0_phase2 : c1990 ? write_point0_phase2 : c1991 ? write_point0_phase2 : c1992 ? write_point0_phase2 : c1993 ? write_point0_phase2 : c1994 ? write_point0_phase2 : c1995 ? write_point0_phase2 : c1996 ? write_point0_phase2 : ((c2055 || c2091) || c2090) ? write_point0_phase2 : c1998 ? write_point0_phase2 : c1999 ? write_point0_phase2 : c2000 ? write_point0_phase2 : c2001 ? write_point0_phase2 : (c2199 || c2198) ? write_point0_phase2 : (c2002 && !c927) ? write_point0_phase2 : c1972 ? write_point0_phase2 : 'bz; */
            /* zero_pop_return0_ip6 <= (c1971 && c889) ? zero_pop_return0_ip2 : ((c2004 || c2005) || c2006) ? zero_pop_return0_ip2 : c1974 ? zero_pop_return0_ip2 : c1975 ? zero_pop_return0_ip2 : c1976 ? zero_pop_return0_ip2 : c1977 ? zero_pop_return0_ip2 : c1978 ? zero_pop_return0_ip2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? zero_pop_return0_ip2 : (((c2019 || c2017) || c2018) || c2016) ? zero_pop_return0_ip2 : c1981 ? zero_pop_return0_ip2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? zero_pop_return0_ip2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? zero_pop_return0_ip2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? zero_pop_return0_ip2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? zero_pop_return0_ip2 : (((c2038 || c2040) || c2037) || c2039) ? zero_pop_return0_ip2 : (c2041 || c2042) ? zero_pop_return0_ip2 : c1988 ? zero_pop_return0_ip2 : c1989 ? zero_pop_return0_ip2 : c1990 ? zero_pop_return0_ip2 : c1991 ? zero_pop_return0_ip2 : c1992 ? zero_pop_return0_ip2 : c1993 ? zero_pop_return0_ip2 : c1994 ? zero_pop_return0_ip2 : c1995 ? zero_pop_return0_ip2 : c1996 ? zero_pop_return0_ip2 : ((c2055 || c2091) || c2090) ? zero_pop_return0_ip5 : c1998 ? zero_pop_return0_ip2 : c1999 ? zero_pop_return0_ip2 : c2000 ? zero_pop_return0_ip2 : c2001 ? zero_pop_return0_ip2 : (c2199 || c2198) ? zero_pop_return0_ip2 : (c2002 && !c927) ? zero_pop_return0_ip2 : c1972 ? zero_pop_return0_ip2 : 'bz; */
            /* zero_pop_return0_phase6 <= (c1971 && c889) ? zero_pop_return0_phase2 : ((c2004 || c2005) || c2006) ? zero_pop_return0_phase2 : c1974 ? zero_pop_return0_phase2 : c1975 ? zero_pop_return0_phase2 : c1976 ? zero_pop_return0_phase2 : c1977 ? zero_pop_return0_phase2 : c1978 ? zero_pop_return0_phase2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? zero_pop_return0_phase2 : (((c2019 || c2017) || c2018) || c2016) ? zero_pop_return0_phase2 : c1981 ? zero_pop_return0_phase2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? zero_pop_return0_phase2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? zero_pop_return0_phase2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? zero_pop_return0_phase2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? zero_pop_return0_phase2 : (((c2038 || c2040) || c2037) || c2039) ? zero_pop_return0_phase2 : (c2041 || c2042) ? zero_pop_return0_phase2 : c1988 ? zero_pop_return0_phase2 : c1989 ? zero_pop_return0_phase2 : c1990 ? zero_pop_return0_phase2 : c1991 ? zero_pop_return0_phase2 : c1992 ? zero_pop_return0_phase2 : c1993 ? zero_pop_return0_phase2 : c1994 ? zero_pop_return0_phase2 : c1995 ? zero_pop_return0_phase2 : c1996 ? zero_pop_return0_phase2 : ((c2055 || c2091) || c2090) ? zero_pop_return0_phase5 : c1998 ? zero_pop_return0_phase2 : c1999 ? zero_pop_return0_phase2 : c2000 ? zero_pop_return0_phase2 : c2001 ? zero_pop_return0_phase2 : (c2199 || c2198) ? zero_pop_return0_phase2 : (c2002 && !c927) ? zero_pop_return0_phase2 : c1972 ? zero_pop_return0_phase2 : 'bz; */
            /* c920 <= (wr_flag4 != 0); */
            /* c2200 <= (c886 && c920); */
            retro_main_state <= retro_main_L1_b178_S1;
          end else if (c1041) begin
            /* c879_inl13 <= (lit0_phase2 == 0); */
            /* c880_inl13 <= (lit0_phase2 == 1); */
            /* c1036_inl13 <= (!c879_inl13 && c880_inl13); */
            /* c1037_inl13 <= (!c879_inl13 && !c880_inl13); */
            /* c3339 <= (c3337 && c1041); */
            /* c1973 <= (c1971 && c1041); */
            if (c879_inl13) begin
              /* lit0_ip3 <= (ip2 + 1); */
              /* c3369 <= (c3339 && c879_inl13); */
              /* c2004 <= (c1973 && c879_inl13); */
              retro_main_state <= retro_main_L1_exit219_S0;
            end else if (c1036_inl13) begin
              /* c3370 <= (c3339 && c1036_inl13); */
              /* c2005 <= (c1973 && c1036_inl13); */
              retro_main_state <= retro_main_L1_exit219_S0;
            end else if (c1037_inl13) begin
              /* c881_inl13 <= (lit0_phase2 == 2); */
              /* stack0_pos3 <= (stack0_pos2 + 1); */
              if (!(lit0_phase2 === 2)) begin
                $display("ASSERTION FAILED (lit0_phase2 === 2)"); $finish;
              end
              /* c3371 <= (c3339 && c1037_inl13); */
              /* c2006 <= (c1973 && c1037_inl13); */
              retro_main_state <= retro_main_L1_ifelse221_S3;
            end
          end else if (c1042) begin
            _stack_addr <= t839_inl14;
            _stack_we <= 1;
            _stack_req <= 1;
            _stack_d <= stack0_second2;
            /* t839_inl14 <= (stack0_pos2 - 2); */
            /* stack0_pos5 <= (stack0_pos2 + 1); */
            /* c3340 <= (c3337 && c1042); */
            /* c1974 <= (c1971 && c1042); */
            retro_main_state <= retro_main_L1_ifthen20_S1;
          end else if (c1043) begin
            _stack_addr <= t842_inl18;
            _stack_we <= 0;
            _stack_req <= 1;
            /* stack0_pos6 <= (stack0_pos2 - 1); */
            /* t842_inl18 <= (stack0_pos6 - 2); */
            /* c3341 <= (c3337 && c1043); */
            /* c1975 <= (c1971 && c1043); */
            retro_main_state <= retro_main_L1_ifthen24_S1;
          end else if (c1044) begin
            /* c3342 <= (c3337 && c1044); */
            /* c1976 <= (c1971 && c1044); */
            retro_main_state <= retro_main_L1_b178_S0;
          end else if (c1045) begin
            _stack_addr <= t842_inl19;
            _stack_we <= 0;
            _stack_req <= 1;
            _address_addr <= t839_inl15;
            _address_we <= 1;
            _address_req <= 1;
            _address_d <= address0_second2;
            /* stack0_pos7 <= (stack0_pos2 - 1); */
            /* t839_inl15 <= (address0_pos2 - 2); */
            /* address0_pos3 <= (address0_pos2 + 1); */
            /* t842_inl19 <= (stack0_pos7 - 2); */
            /* c3343 <= (c3337 && c1045); */
            /* c1977 <= (c1971 && c1045); */
            retro_main_state <= retro_main_L1_ifthen32_S1;
          end else if (c1046) begin
            _address_addr <= t842_inl20;
            _address_we <= 0;
            _address_req <= 1;
            _stack_addr <= t839_inl16;
            _stack_we <= 1;
            _stack_req <= 1;
            _stack_d <= stack0_second2;
            /* address0_pos4 <= (address0_pos2 - 1); */
            /* t839_inl16 <= (stack0_pos2 - 2); */
            /* stack0_pos8 <= (stack0_pos2 + 1); */
            /* t842_inl20 <= (address0_pos4 - 2); */
            /* c3344 <= (c3337 && c1046); */
            /* c1978 <= (c1971 && c1046); */
            retro_main_state <= retro_main_L1_ifthen36_S1;
          end else if (c1047) begin
            /* c872_inl33 <= (loop0_phase2 == 0); */
            /* c873_inl33 <= (loop0_phase2 == 1); */
            /* c874_inl33 <= (loop0_phase2 == 2); */
            /* c1033_inl33 <= (!c872_inl33 && c873_inl33); */
            /* c1034_inl33 <= ((!c872_inl33 && !c873_inl33) && c874_inl33); */
            /* c1035_inl33 <= ((!c872_inl33 && !c873_inl33) && !c874_inl33); */
            /* c3345 <= (c3337 && c1047); */
            /* c1979 <= (c1971 && c1047); */
            if (c872_inl33) begin
              /* loop0_ip3 <= (ip2 + 1); */
              /* c3372 <= (c3345 && c872_inl33); */
              /* c2012 <= (c1979 && c872_inl33); */
              retro_main_state <= retro_main_L1_ifthen304_S3;
            end else if (c1033_inl33) begin
              /* c3373 <= (c3345 && c1033_inl33); */
              /* c2013 <= (c1979 && c1033_inl33); */
              retro_main_state <= retro_main_L1_exit310_S0;
            end else if (c1034_inl33) begin
              /* c3374 <= (c3345 && c1034_inl33); */
              /* c2014 <= (c1979 && c1034_inl33); */
              retro_main_state <= retro_main_L1_ifthen317_S7;
            end else if (c1035_inl33) begin
              /* c878_inl33 <= (loop0_phase2 == 3); */
              if (!(loop0_phase2 === 3)) begin
                $display("ASSERTION FAILED (loop0_phase2 === 3)"); $finish;
              end
              /* c3375 <= (c3345 && c1035_inl33); */
              /* c2015 <= (c1979 && c1035_inl33); */
              retro_main_state <= retro_main_L1_exit310_S0;
            end
          end else if (c1048) begin
            /* c882_inl34 <= (jump0_phase2 == 0); */
            /* c883_inl34 <= (jump0_phase2 == 1); */
            /* c884_inl34 <= (jump0_phase2 == 2); */
            /* jump0_ip3 <= (ip2 + 1); */
            /* c885_inl34 <= (jump0_phase2 == 3); */
            /* c1038_inl34 <= (!c882_inl34 && c883_inl34); */
            /* c1039_inl34 <= ((!c882_inl34 && !c883_inl34) && c884_inl34); */
            /* c1040_inl34 <= ((!c882_inl34 && !c883_inl34) && !c884_inl34); */
            /* c3346 <= (c3337 && c1048); */
            /* c1980 <= (c1971 && c1048); */
            /* c2016 <= (c1980 && c882_inl34); */
            /* c2017 <= (c1980 && c1038_inl34); */
            /* c2018 <= (c1980 && c1039_inl34); */
            /* c2019 <= (c1980 && c1040_inl34); */
            retro_main_state <= retro_main_L1_ifthen44_S1;
          end else if (c1049) begin
            /* c3347 <= (c3337 && c1049); */
            /* c1981 <= (c1971 && c1049); */
            retro_main_state <= retro_main_L1_ifthen48_S1;
          end else if (c1050) begin
            /* c867_inl35 <= (jump_ge0_phase2 == 0); */
            /* c868_inl35 <= (jump_ge0_phase2 == 1); */
            /* c869_inl35 <= (jump_ge0_phase2 == 2); */
            /* c1030_inl35 <= (!c867_inl35 && c868_inl35); */
            /* c1031_inl35 <= ((!c867_inl35 && !c868_inl35) && c869_inl35); */
            /* c1032_inl35 <= ((!c867_inl35 && !c868_inl35) && !c869_inl35); */
            /* c3348 <= (c3337 && c1050); */
            /* c1982 <= (c1971 && c1050); */
            if (c867_inl35) begin
              /* c3377 <= (c3348 && c867_inl35); */
              /* c2021 <= (c1982 && c867_inl35); */
              retro_main_state <= retro_main_L1_ifthen328_S1;
            end else if (c1030_inl35) begin
              /* c870_inl35 <= (stack0_top2 > jump_ge0_a2); */
              /* c3378 <= (c3348 && c1030_inl35); */
              /* c2022 <= (c1982 && c1030_inl35); */
              /* c2126 <= (c2022 && c870_inl35); */
              /* c2127 <= (c2022 && !c870_inl35); */
              retro_main_state <= retro_main_L1_ifthen334_S4;
            end else if (c1031_inl35) begin
              /* c3379 <= (c3348 && c1031_inl35); */
              /* c2023 <= (c1982 && c1031_inl35); */
              retro_main_state <= retro_main_L1_ifthen341_S7;
            end else if (c1032_inl35) begin
              /* c871_inl35 <= (jump_ge0_phase2 == 3); */
              if (!(jump_ge0_phase2 === 3)) begin
                $display("ASSERTION FAILED (jump_ge0_phase2 === 3)"); $finish;
              end
              /* c3380 <= (c3348 && c1032_inl35); */
              /* c2024 <= (c1982 && c1032_inl35); */
              retro_main_state <= retro_main_L1_exit333_S0;
            end
          end else if (c1051) begin
            /* c862_inl36 <= (jump_le0_phase2 == 0); */
            /* c863_inl36 <= (jump_le0_phase2 == 1); */
            /* c864_inl36 <= (jump_le0_phase2 == 2); */
            /* c1027_inl36 <= (!c862_inl36 && c863_inl36); */
            /* c1028_inl36 <= ((!c862_inl36 && !c863_inl36) && c864_inl36); */
            /* c1029_inl36 <= ((!c862_inl36 && !c863_inl36) && !c864_inl36); */
            /* c3349 <= (c3337 && c1051); */
            /* c1983 <= (c1971 && c1051); */
            if (c862_inl36) begin
              /* c3381 <= (c3349 && c862_inl36); */
              /* c2025 <= (c1983 && c862_inl36); */
              retro_main_state <= retro_main_L1_ifthen345_S1;
            end else if (c1027_inl36) begin
              /* c865_inl36 <= (stack0_top2 < jump_le0_a2); */
              /* c3382 <= (c3349 && c1027_inl36); */
              /* c2026 <= (c1983 && c1027_inl36); */
              /* c2128 <= (c2026 && c865_inl36); */
              /* c2129 <= (c2026 && !c865_inl36); */
              retro_main_state <= retro_main_L1_ifthen351_S4;
            end else if (c1028_inl36) begin
              /* c3383 <= (c3349 && c1028_inl36); */
              /* c2027 <= (c1983 && c1028_inl36); */
              retro_main_state <= retro_main_L1_ifthen358_S7;
            end else if (c1029_inl36) begin
              /* c866_inl36 <= (jump_le0_phase2 == 3); */
              if (!(jump_le0_phase2 === 3)) begin
                $display("ASSERTION FAILED (jump_le0_phase2 === 3)"); $finish;
              end
              /* c3384 <= (c3349 && c1029_inl36); */
              /* c2028 <= (c1983 && c1029_inl36); */
              retro_main_state <= retro_main_L1_exit350_S0;
            end
          end else if (c1052) begin
            /* c857_inl37 <= (jump_ne0_phase2 == 0); */
            /* c858_inl37 <= (jump_ne0_phase2 == 1); */
            /* c859_inl37 <= (jump_ne0_phase2 == 2); */
            /* c1024_inl37 <= (!c857_inl37 && c858_inl37); */
            /* c1025_inl37 <= ((!c857_inl37 && !c858_inl37) && c859_inl37); */
            /* c1026_inl37 <= ((!c857_inl37 && !c858_inl37) && !c859_inl37); */
            /* c3350 <= (c3337 && c1052); */
            /* c1984 <= (c1971 && c1052); */
            if (c857_inl37) begin
              /* c3385 <= (c3350 && c857_inl37); */
              /* c2029 <= (c1984 && c857_inl37); */
              retro_main_state <= retro_main_L1_ifthen362_S1;
            end else if (c1024_inl37) begin
              /* c860_inl37 <= (stack0_top2 != jump_ne0_a2); */
              /* c3386 <= (c3350 && c1024_inl37); */
              /* c2030 <= (c1984 && c1024_inl37); */
              /* c2130 <= (c2030 && c860_inl37); */
              /* c2131 <= (c2030 && !c860_inl37); */
              retro_main_state <= retro_main_L1_ifthen368_S4;
            end else if (c1025_inl37) begin
              /* c3387 <= (c3350 && c1025_inl37); */
              /* c2031 <= (c1984 && c1025_inl37); */
              retro_main_state <= retro_main_L1_ifthen375_S7;
            end else if (c1026_inl37) begin
              /* c861_inl37 <= (jump_ne0_phase2 == 3); */
              if (!(jump_ne0_phase2 === 3)) begin
                $display("ASSERTION FAILED (jump_ne0_phase2 === 3)"); $finish;
              end
              /* c3388 <= (c3350 && c1026_inl37); */
              /* c2032 <= (c1984 && c1026_inl37); */
              retro_main_state <= retro_main_L1_exit367_S0;
            end
          end else if (c1053) begin
            /* c852_inl38 <= (jump_eq0_phase2 == 0); */
            /* c853_inl38 <= (jump_eq0_phase2 == 1); */
            /* c854_inl38 <= (jump_eq0_phase2 == 2); */
            /* c1021_inl38 <= (!c852_inl38 && c853_inl38); */
            /* c1022_inl38 <= ((!c852_inl38 && !c853_inl38) && c854_inl38); */
            /* c1023_inl38 <= ((!c852_inl38 && !c853_inl38) && !c854_inl38); */
            /* c3351 <= (c3337 && c1053); */
            /* c1985 <= (c1971 && c1053); */
            if (c852_inl38) begin
              /* c3389 <= (c3351 && c852_inl38); */
              /* c2033 <= (c1985 && c852_inl38); */
              retro_main_state <= retro_main_L1_ifthen379_S1;
            end else if (c1021_inl38) begin
              /* c855_inl38 <= (stack0_top2 == jump_eq0_a2); */
              /* c3390 <= (c3351 && c1021_inl38); */
              /* c2034 <= (c1985 && c1021_inl38); */
              /* c2132 <= (c2034 && c855_inl38); */
              /* c2133 <= (c2034 && !c855_inl38); */
              retro_main_state <= retro_main_L1_ifthen385_S5;
            end else if (c1022_inl38) begin
              /* c3391 <= (c3351 && c1022_inl38); */
              /* c2035 <= (c1985 && c1022_inl38); */
              retro_main_state <= retro_main_L1_ifthen392_S7;
            end else if (c1023_inl38) begin
              /* c856_inl38 <= (jump_eq0_phase2 == 3); */
              if (!(jump_eq0_phase2 === 3)) begin
                $display("ASSERTION FAILED (jump_eq0_phase2 === 3)"); $finish;
              end
              /* c3392 <= (c3351 && c1023_inl38); */
              /* c2036 <= (c1985 && c1023_inl38); */
              retro_main_state <= retro_main_L1_exit384_S0;
            end
          end else if (c1054) begin
            /* c848_inl39 <= (point0_phase2 == 0); */
            /* c849_inl39 <= (point0_phase2 == 1); */
            /* c850_inl39 <= (point0_phase2 == 2); */
            /* c1018_inl39 <= (!c848_inl39 && c849_inl39); */
            /* c1019_inl39 <= ((!c848_inl39 && !c849_inl39) && c850_inl39); */
            /* c1020_inl39 <= ((!c848_inl39 && !c849_inl39) && !c850_inl39); */
            /* c3352 <= (c3337 && c1054); */
            /* c1986 <= (c1971 && c1054); */
            if (c848_inl39) begin
              /* c3393 <= (c3352 && c848_inl39); */
              /* c2037 <= (c1986 && c848_inl39); */
              retro_main_state <= retro_main_L1_exit397_S0;
            end else if (c1018_inl39) begin
              /* c3394 <= (c3352 && c1018_inl39); */
              /* c2038 <= (c1986 && c1018_inl39); */
              retro_main_state <= retro_main_L1_exit397_S0;
            end else if (c1019_inl39) begin
              /* c3395 <= (c3352 && c1019_inl39); */
              /* c2039 <= (c1986 && c1019_inl39); */
              retro_main_state <= retro_main_L1_exit397_S0;
            end else if (c1020_inl39) begin
              /* c851_inl39 <= (point0_phase2 == 3); */
              if (!(point0_phase2 === 3)) begin
                $display("ASSERTION FAILED (point0_phase2 === 3)"); $finish;
              end
              /* c3396 <= (c3352 && c1020_inl39); */
              /* c2040 <= (c1986 && c1020_inl39); */
              retro_main_state <= retro_main_L1_exit397_S0;
            end
          end else if (c1055) begin
            /* c843_inl40 <= (write_point0_phase2 == 0); */
            /* c3353 <= (c3337 && c1055); */
            /* c1987 <= (c1971 && c1055); */
            if (c843_inl40) begin
              /* c3397 <= (c3353 && c843_inl40); */
              /* c2041 <= (c1987 && c843_inl40); */
              retro_main_state <= retro_main_L1_ifthen407_S5;
            end else begin
              /* c844_inl40 <= (write_point0_phase2 == 1); */
              if (!(write_point0_phase2 === 1)) begin
                $display("ASSERTION FAILED (write_point0_phase2 === 1)"); $finish;
              end
              /* c3398 <= (c3353 && !c843_inl40); */
              /* c2042 <= (c1987 && !c843_inl40); */
              retro_main_state <= retro_main_L1_ifelse413_S5;
            end
          end else if (c1056) begin
            /* stack0_top31 <= (stack0_second2 + stack0_top2); */
            /* c3354 <= (c3337 && c1056); */
            /* c1988 <= (c1971 && c1056); */
            retro_main_state <= retro_main_L1_ifthen81_S1;
          end else if (c1057) begin
            /* c3355 <= (c3337 && c1057); */
            /* c1989 <= (c1971 && c1057); */
            retro_main_state <= retro_main_L1_ifthen85_S1;
          end else if (c1058) begin
            /* stack0_top35 <= (stack0_second2 * stack0_top2); */
            /* c3356 <= (c3337 && c1058); */
            /* c1990 <= (c1971 && c1058); */
            retro_main_state <= retro_main_L1_ifthen89_S1;
          end else if (c1059) begin
            /* c1005_inl1_inl52 <= (stack0_second2 < 0); */
            /* c1005_inl2_inl52 <= (stack0_top2 < 0); */
            /* c996_inl52 <= (stack0_second2 < 0); */
            /* c997_inl52 <= (stack0_top2 < 0); */
            /* c999_inl52 <= (stack0_second2 > 0); */
            /* c1000_inl52 <= (stack0_top2 < 0); */
            /* c1002_inl52 <= (stack0_second2 < 0); */
            /* c1003_inl52 <= (stack0_top2 > 0); */
            /* t1006_inl1_inl52 <= c1005_inl1_inl52 ? -stack0_second2 : stack0_second2; */
            /* t1006_inl2_inl52 <= c1005_inl2_inl52 ? -stack0_top2 : stack0_top2; */
            /* c998_inl52 <= (c996_inl52 && c997_inl52); */
            /* c1001_inl52 <= (c999_inl52 && c1000_inl52); */
            /* c1004_inl52 <= (c1002_inl52 && c1003_inl52); */
            /* q_inl522 <= (t1006_inl1_inl52 / t1006_inl2_inl52); */
            /* r_inl522 <= (t1006_inl1_inl52 % t1006_inl2_inl52); */
            /* c1094_inl52 <= (!c998_inl52 && c1001_inl52); */
            /* c1095_inl52 <= ((!c998_inl52 && !c1001_inl52) && c1004_inl52); */
            /* c1096_inl52 <= ((!c998_inl52 && !c1001_inl52) && !c1004_inl52); */
            /* r_inl523 <= (r_inl522 * -1); */
            /* q_inl523 <= (q_inl522 * -1); */
            /* r_inl524 <= (r_inl522 * -1); */
            /* q_inl524 <= (q_inl522 * -1); */
            /* c3357 <= (c3337 && c1059); */
            /* c1991 <= (c1971 && c1059); */
            /* c2046 <= (c1991 && c998_inl52); */
            /* c2047 <= (c1991 && c1094_inl52); */
            /* c2048 <= (c1991 && c1095_inl52); */
            /* q_inl525 <= c2046 ? q_inl522 : c2047 ? q_inl523 : c2048 ? q_inl524 : (c1991 && c1096_inl52) ? q_inl522 : 'bz; */
            /* r_inl525 <= c2046 ? r_inl523 : c2047 ? r_inl522 : c2048 ? r_inl524 : (c1991 && c1096_inl52) ? r_inl522 : 'bz; */
            array1007_inl52[0] <= q_inl525;
            array1007_inl52[1] <= r_inl525;
            retro_main_state <= retro_main_L1_ifthen93_S2;
          end else if (c1060) begin
            /* stack0_top38 <= (stack0_second2 & stack0_top2); */
            /* c3358 <= (c3337 && c1060); */
            /* c1992 <= (c1971 && c1060); */
            retro_main_state <= retro_main_L1_ifthen97_S2;
          end else if (c1061) begin
            /* stack0_top40 <= (stack0_second2 | stack0_top2); */
            /* c3359 <= (c3337 && c1061); */
            /* c1993 <= (c1971 && c1061); */
            retro_main_state <= retro_main_L1_ifthen101_S2;
          end else if (c1062) begin
            /* stack0_top42 <= (stack0_second2 ^ stack0_top2); */
            /* c3360 <= (c3337 && c1062); */
            /* c1994 <= (c1971 && c1062); */
            retro_main_state <= retro_main_L1_ifthen105_S2;
          end else if (c1063) begin
            /* stack0_top44 <= (stack0_second2 << stack0_top2); */
            /* c3361 <= (c3337 && c1063); */
            /* c1995 <= (c1971 && c1063); */
            retro_main_state <= retro_main_L1_ifthen109_S2;
          end else if (c1064) begin
            /* stack0_top46 <= (stack0_second2 >>> stack0_top2); */
            /* c3362 <= (c3337 && c1064); */
            /* c1996 <= (c1971 && c1064); */
            retro_main_state <= retro_main_L1_ifthen113_S2;
          end else if (c1065) begin
            /* c845_inl54 <= (zero_pop_return0_phase2 == 0); */
            /* c3363 <= (c3337 && c1065); */
            /* c1997 <= (c1971 && c1065); */
            if (c845_inl54) begin
              /* c846_inl54 <= (stack0_top2 == 0); */
              /* c3399 <= (c3363 && c845_inl54); */
              /* c2054 <= (c1997 && c845_inl54); */
              if (c846_inl54) begin
                /* c3405 <= (c3399 && c846_inl54); */
                /* c2090 <= (c2054 && c846_inl54); */
                retro_main_state <= retro_main_L1_ifthen479_S6;
              end else begin
                /* c3406 <= (c3399 && !c846_inl54); */
                /* c2091 <= (c2054 && !c846_inl54); */
                retro_main_state <= retro_main_L1_exit488_S0;
              end
            end else begin
              /* c847_inl54 <= (zero_pop_return0_phase2 == 1); */
              if (!(zero_pop_return0_phase2 === 1)) begin
                $display("ASSERTION FAILED (zero_pop_return0_phase2 === 1)"); $finish;
              end
              /* c3400 <= (c3363 && !c845_inl54); */
              /* c2055 <= (c1997 && !c845_inl54); */
              retro_main_state <= retro_main_L1_exit488_S0;
            end
          end else if (c1066) begin
            /* stack0_top49 <= (stack0_top2 + 1); */
            /* c3364 <= (c3337 && c1066); */
            /* c1998 <= (c1971 && c1066); */
            retro_main_state <= retro_main_L1_b178_S0;
          end else if (c1067) begin
            /* c3365 <= (c3337 && c1067); */
            /* c1999 <= (c1971 && c1067); */
            retro_main_state <= retro_main_L1_ifthen125_S3;
          end else if (c1068) begin
            stack0_top51 <= array1010[stack0_top2];
            array1010[stack0_top2] <= 0;
            /* c3366 <= (c3337 && c1068); */
            /* c2000 <= (c1971 && c1068); */
            retro_main_state <= retro_main_L1_b178_S0;
          end else if (c1069) begin
            array1010[stack0_top2] <= stack0_second2;
            /* c3367 <= (c3337 && c1069); */
            /* c2001 <= (c1971 && c1069); */
            retro_main_state <= retro_main_L1_ifthen133_S3;
          end else if (c1070) begin
            t926 <= array1010[0];
            /* c3368 <= (c3337 && c1070); */
            /* c2002 <= (c1971 && c1070); */
            retro_main_state <= retro_main_L1_ifthen137_S1;
          end else if (c1071) begin
            retro_main_valid <= 1;
            if (retro_main_accept == 1) begin
              retro_main_state <= retro_main_b1_INIT;
            end
          end
        end else begin
          _address_addr <= t839_inl17;
          _address_we <= 1;
          _address_req <= 1;
          _address_d <= address0_second2;
          memory_addr <= ip2;
          memory_we <= 0;
          memory_req <= 1;
          /* t839_inl17 <= (address0_pos2 - 2); */
          /* address0_pos8 <= (address0_pos2 + 1); */
          /* c3338 <= (c886 && !c888); */
          /* c1972 <= (c886 && !c888); */
          retro_main_state <= retro_main_L1_ifelse177_S1;
        end
      end
      retro_main_L1_ifelse177_S1: begin
        _address_req <= 0;
        /*wait for output of memory*/
        retro_main_state <= retro_main_L1_ifelse177_S2;
      end
      retro_main_L1_ifelse177_S2: begin
        t928 <= memory_q;
        memory_req <= 0;
        retro_main_state <= retro_main_L1_ifelse177_S3;
      end
      retro_main_L1_ifelse177_S3: begin
        /* ip15 <= (t928 - 1); */
        retro_main_state <= retro_main_L1_b178_S0;
      end
      retro_main_L1_ifthen20_S1: begin
        _stack_req <= 0;
        retro_main_state <= retro_main_L1_b178_S0;
      end
      retro_main_L1_ifthen24_S1: begin
        /*wait for output of _stack*/
        retro_main_state <= retro_main_L1_ifthen24_S2;
      end
      retro_main_L1_ifthen24_S2: begin
        stack0_second6 <= _stack_q;
        _stack_req <= 0;
        retro_main_state <= retro_main_L1_b178_S0;
      end
      retro_main_L1_ifthen32_S1: begin
        /*wait for output of _stack*/
        _address_req <= 0;
        retro_main_state <= retro_main_L1_ifthen32_S2;
      end
      retro_main_L1_ifthen32_S2: begin
        stack0_second8 <= _stack_q;
        _stack_req <= 0;
        retro_main_state <= retro_main_L1_b178_S0;
      end
      retro_main_L1_ifthen36_S1: begin
        /*wait for output of _address*/
        _stack_req <= 0;
        retro_main_state <= retro_main_L1_ifthen36_S2;
      end
      retro_main_L1_ifthen36_S2: begin
        address0_second4 <= _address_q;
        _address_req <= 0;
        retro_main_state <= retro_main_L1_b178_S0;
      end
      retro_main_L1_ifthen44_S1: begin
        /* jump0_ip4 <= (mem_data - 1); */
        if (c882_inl34) begin
          /* c3404 <= (((c3346 && c882_inl34) || (c3346 && c1038_inl34)) || (c3346 && c1039_inl34)); */
          /* exec_result346 <= c2016 ? 0 : c2017 ? 0 : c2018 ? 0 : c2019 ? 1 : 'bz; */
          /* jump0_ip5 <= c2016 ? jump0_ip3 : c2017 ? jump0_ip2 : c2018 ? jump0_ip4 : c2019 ? jump0_ip2 : 'bz; */
          /* jump0_phase7 <= c2016 ? 1 : c2017 ? 2 : c2018 ? 3 : c2019 ? 0 : 'bz; */
          retro_main_state <= retro_main_L1_b178_S0;
        end else if (c1038_inl34) begin
          /* c3404 <= (((c3346 && c882_inl34) || (c3346 && c1038_inl34)) || (c3346 && c1039_inl34)); */
          /* exec_result346 <= c2016 ? 0 : c2017 ? 0 : c2018 ? 0 : c2019 ? 1 : 'bz; */
          /* jump0_ip5 <= c2016 ? jump0_ip3 : c2017 ? jump0_ip2 : c2018 ? jump0_ip4 : c2019 ? jump0_ip2 : 'bz; */
          /* jump0_phase7 <= c2016 ? 1 : c2017 ? 2 : c2018 ? 3 : c2019 ? 0 : 'bz; */
          retro_main_state <= retro_main_L1_b178_S0;
        end else if (c1039_inl34) begin
          /* c3404 <= (((c3346 && c882_inl34) || (c3346 && c1038_inl34)) || (c3346 && c1039_inl34)); */
          /* exec_result346 <= c2016 ? 0 : c2017 ? 0 : c2018 ? 0 : c2019 ? 1 : 'bz; */
          /* jump0_ip5 <= c2016 ? jump0_ip3 : c2017 ? jump0_ip2 : c2018 ? jump0_ip4 : c2019 ? jump0_ip2 : 'bz; */
          /* jump0_phase7 <= c2016 ? 1 : c2017 ? 2 : c2018 ? 3 : c2019 ? 0 : 'bz; */
          retro_main_state <= retro_main_L1_b178_S0;
        end else if (c1040_inl34) begin
          if (!(jump0_phase2 === 3)) begin
            $display("ASSERTION FAILED (jump0_phase2 === 3)"); $finish;
          end
          /* c3376 <= (c3346 && c1040_inl34); */
          retro_main_state <= retro_main_L1_exit322_S0;
        end
      end
      retro_main_L1_ifthen48_S1: begin
        _address_addr <= t842_inl21;
        _address_we <= 0;
        _address_req <= 1;
        /* address0_pos5 <= (address0_pos2 - 1); */
        /* t842_inl21 <= (address0_pos5 - 2); */
        retro_main_state <= retro_main_L1_ifthen48_S2;
      end
      retro_main_L1_ifthen48_S2: begin
        /*wait for output of _address*/
        retro_main_state <= retro_main_L1_ifthen48_S3;
      end
      retro_main_L1_ifthen48_S3: begin
        address0_second5 <= _address_q;
        _address_req <= 0;
        retro_main_state <= retro_main_L1_b178_S0;
      end
      retro_main_L1_ifthen81_S1: begin
        _stack_addr <= t842_inl22;
        _stack_we <= 0;
        _stack_req <= 1;
        /* stack0_pos26 <= (stack0_pos2 - 1); */
        /* t842_inl22 <= (stack0_pos26 - 2); */
        retro_main_state <= retro_main_L1_ifthen81_S2;
      end
      retro_main_L1_ifthen81_S2: begin
        /*wait for output of _stack*/
        retro_main_state <= retro_main_L1_ifthen81_S3;
      end
      retro_main_L1_ifthen81_S3: begin
        stack0_second27 <= _stack_q;
        _stack_req <= 0;
        retro_main_state <= retro_main_L1_b178_S0;
      end
      retro_main_L1_ifthen85_S1: begin
        _stack_addr <= t842_inl23;
        _stack_we <= 0;
        _stack_req <= 1;
        /* stack0_pos27 <= (stack0_pos2 - 1); */
        /* stack0_top33 <= (stack0_second2 - stack0_top2); */
        /* t842_inl23 <= (stack0_pos27 - 2); */
        retro_main_state <= retro_main_L1_ifthen85_S2;
      end
      retro_main_L1_ifthen85_S2: begin
        /*wait for output of _stack*/
        retro_main_state <= retro_main_L1_ifthen85_S3;
      end
      retro_main_L1_ifthen85_S3: begin
        stack0_second28 <= _stack_q;
        _stack_req <= 0;
        retro_main_state <= retro_main_L1_b178_S0;
      end
      retro_main_L1_ifthen89_S1: begin
        _stack_addr <= t842_inl24;
        _stack_we <= 0;
        _stack_req <= 1;
        /* stack0_pos28 <= (stack0_pos2 - 1); */
        /* t842_inl24 <= (stack0_pos28 - 2); */
        retro_main_state <= retro_main_L1_ifthen89_S2;
      end
      retro_main_L1_ifthen89_S2: begin
        /*wait for output of _stack*/
        retro_main_state <= retro_main_L1_ifthen89_S3;
      end
      retro_main_L1_ifthen89_S3: begin
        stack0_second29 <= _stack_q;
        _stack_req <= 0;
        retro_main_state <= retro_main_L1_b178_S0;
      end
      retro_main_L1_ifthen93_S2: begin
        /* stack0_top36 <= retro_divmod_result522[0]; */
        /* stack0_second30 <= retro_divmod_result522[1]; */
        retro_main_state <= retro_main_L1_b178_S0;
      end
      retro_main_L1_ifthen97_S2: begin
        _stack_addr <= t842_inl25;
        _stack_we <= 0;
        _stack_req <= 1;
        /* stack0_pos29 <= (stack0_pos2 - 1); */
        /* t842_inl25 <= (stack0_pos29 - 2); */
        retro_main_state <= retro_main_L1_ifthen97_S3;
      end
      retro_main_L1_ifthen97_S3: begin
        /*wait for output of _stack*/
        retro_main_state <= retro_main_L1_ifthen97_S4;
      end
      retro_main_L1_ifthen97_S4: begin
        stack0_second31 <= _stack_q;
        _stack_req <= 0;
        retro_main_state <= retro_main_L1_b178_S0;
      end
      retro_main_L1_ifthen101_S2: begin
        _stack_addr <= t842_inl26;
        _stack_we <= 0;
        _stack_req <= 1;
        /* stack0_pos30 <= (stack0_pos2 - 1); */
        /* t842_inl26 <= (stack0_pos30 - 2); */
        retro_main_state <= retro_main_L1_ifthen101_S3;
      end
      retro_main_L1_ifthen101_S3: begin
        /*wait for output of _stack*/
        retro_main_state <= retro_main_L1_ifthen101_S4;
      end
      retro_main_L1_ifthen101_S4: begin
        stack0_second32 <= _stack_q;
        _stack_req <= 0;
        retro_main_state <= retro_main_L1_b178_S0;
      end
      retro_main_L1_ifthen105_S2: begin
        _stack_addr <= t842_inl27;
        _stack_we <= 0;
        _stack_req <= 1;
        /* stack0_pos31 <= (stack0_pos2 - 1); */
        /* t842_inl27 <= (stack0_pos31 - 2); */
        retro_main_state <= retro_main_L1_ifthen105_S3;
      end
      retro_main_L1_ifthen105_S3: begin
        /*wait for output of _stack*/
        retro_main_state <= retro_main_L1_ifthen105_S4;
      end
      retro_main_L1_ifthen105_S4: begin
        stack0_second33 <= _stack_q;
        _stack_req <= 0;
        retro_main_state <= retro_main_L1_b178_S0;
      end
      retro_main_L1_ifthen109_S2: begin
        _stack_addr <= t842_inl28;
        _stack_we <= 0;
        _stack_req <= 1;
        /* stack0_pos32 <= (stack0_pos2 - 1); */
        /* t842_inl28 <= (stack0_pos32 - 2); */
        retro_main_state <= retro_main_L1_ifthen109_S3;
      end
      retro_main_L1_ifthen109_S3: begin
        /*wait for output of _stack*/
        retro_main_state <= retro_main_L1_ifthen109_S4;
      end
      retro_main_L1_ifthen109_S4: begin
        stack0_second34 <= _stack_q;
        _stack_req <= 0;
        retro_main_state <= retro_main_L1_b178_S0;
      end
      retro_main_L1_ifthen113_S2: begin
        _stack_addr <= t842_inl29;
        _stack_we <= 0;
        _stack_req <= 1;
        /* stack0_pos33 <= (stack0_pos2 - 1); */
        /* t842_inl29 <= (stack0_pos33 - 2); */
        retro_main_state <= retro_main_L1_ifthen113_S3;
      end
      retro_main_L1_ifthen113_S3: begin
        /*wait for output of _stack*/
        retro_main_state <= retro_main_L1_ifthen113_S4;
      end
      retro_main_L1_ifthen113_S4: begin
        stack0_second35 <= _stack_q;
        _stack_req <= 0;
        retro_main_state <= retro_main_L1_b178_S0;
      end
      retro_main_L1_ifthen125_S3: begin
        /* stack0_top50 <= (stack0_top2 - 1); */
        retro_main_state <= retro_main_L1_b178_S0;
      end
      retro_main_L1_ifthen133_S3: begin
        _stack_addr <= t842_inl30;
        _stack_we <= 0;
        _stack_req <= 1;
        /* stack0_pos36 <= (stack0_pos2 - 1); */
        /* t842_inl30 <= (stack0_pos36 - 2); */
        /* stack0_pos37 <= (stack0_pos36 - 1); */
        /* t842_inl31 <= (stack0_pos37 - 2); */
        retro_main_state <= retro_main_L1_ifthen133_S4;
      end
      retro_main_L1_ifthen133_S4: begin
        _stack_addr <= t842_inl31;
        _stack_we <= 0;
        _stack_req <= 1;
        /*wait for output of _stack*/
        retro_main_state <= retro_main_L1_ifthen133_S5;
      end
      retro_main_L1_ifthen133_S5: begin
        /*wait for output of _stack*/
        stack0_second38 <= _stack_q;
        retro_main_state <= retro_main_L1_ifthen133_S6;
      end
      retro_main_L1_ifthen133_S6: begin
        stack0_second39 <= _stack_q;
        _stack_req <= 0;
        retro_main_state <= retro_main_L1_b178_S0;
      end
      retro_main_L1_ifthen137_S1: begin
        /* c927 <= (t926 == 0); */
        if (c927) begin
          array1010[0] <= 1;
          t929_inl55 <= array1010[1];
          /* c3401 <= (c3368 && c927); */
          /* c2060 <= (c2002 && c927); */
          retro_main_state <= retro_main_L1_ifthen140_S1;
        end else begin
          /* address0_pos9 <= (c1971 && c889) ? address0_pos2 : ((c2004 || c2005) || c2006) ? address0_pos2 : c1974 ? address0_pos2 : c1975 ? address0_pos2 : c1976 ? address0_pos2 : c1977 ? address0_pos3 : c1978 ? address0_pos4 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? address0_pos2 : (((c2019 || c2017) || c2018) || c2016) ? address0_pos2 : c1981 ? address0_pos5 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? address0_pos2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? address0_pos2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? address0_pos2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? address0_pos2 : (((c2038 || c2040) || c2037) || c2039) ? address0_pos2 : (c2041 || c2042) ? address0_pos2 : c1988 ? address0_pos2 : c1989 ? address0_pos2 : c1990 ? address0_pos2 : c1991 ? address0_pos2 : c1992 ? address0_pos2 : c1993 ? address0_pos2 : c1994 ? address0_pos2 : c1995 ? address0_pos2 : c1996 ? address0_pos2 : ((c2055 || c2091) || c2090) ? address0_pos7 : c1998 ? address0_pos2 : c1999 ? address0_pos2 : c2000 ? address0_pos2 : c2001 ? address0_pos2 : (c2199 || c2198) ? address0_pos2 : (c2002 && !c927) ? address0_pos2 : c1972 ? address0_pos8 : 'bz; */
          /* address0_second9 <= (c1971 && c889) ? address0_second2 : ((c2004 || c2005) || c2006) ? address0_second2 : c1974 ? address0_second2 : c1975 ? address0_second2 : c1976 ? address0_second2 : c1977 ? address0_top2 : c1978 ? address0_second4 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? address0_second2 : (((c2019 || c2017) || c2018) || c2016) ? address0_second2 : c1981 ? address0_second5 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? address0_second2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? address0_second2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? address0_second2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? address0_second2 : (((c2038 || c2040) || c2037) || c2039) ? address0_second2 : (c2041 || c2042) ? address0_second2 : c1988 ? address0_second2 : c1989 ? address0_second2 : c1990 ? address0_second2 : c1991 ? address0_second2 : c1992 ? address0_second2 : c1993 ? address0_second2 : c1994 ? address0_second2 : c1995 ? address0_second2 : c1996 ? address0_second2 : ((c2055 || c2091) || c2090) ? address0_second7 : c1998 ? address0_second2 : c1999 ? address0_second2 : c2000 ? address0_second2 : c2001 ? address0_second2 : (c2199 || c2198) ? address0_second2 : (c2002 && !c927) ? address0_second2 : c1972 ? address0_top2 : 'bz; */
          /* address0_top9 <= (c1971 && c889) ? address0_top2 : ((c2004 || c2005) || c2006) ? address0_top2 : c1974 ? address0_top2 : c1975 ? address0_top2 : c1976 ? address0_top2 : c1977 ? stack0_top2 : c1978 ? address0_second2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? address0_top2 : (((c2019 || c2017) || c2018) || c2016) ? address0_top2 : c1981 ? address0_second2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? address0_top2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? address0_top2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? address0_top2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? address0_top2 : (((c2038 || c2040) || c2037) || c2039) ? address0_top2 : (c2041 || c2042) ? address0_top2 : c1988 ? address0_top2 : c1989 ? address0_top2 : c1990 ? address0_top2 : c1991 ? address0_top2 : c1992 ? address0_top2 : c1993 ? address0_top2 : c1994 ? address0_top2 : c1995 ? address0_top2 : c1996 ? address0_top2 : ((c2055 || c2091) || c2090) ? address0_top7 : c1998 ? address0_top2 : c1999 ? address0_top2 : c2000 ? address0_top2 : c2001 ? address0_top2 : (c2199 || c2198) ? address0_top2 : (c2002 && !c927) ? address0_top2 : c1972 ? ip2 : 'bz; */
          /* done_flag13 <= (c1971 && c889) ? done_flag2 : ((c2004 || c2005) || c2006) ? exec_result135 : c1974 ? done_flag2 : c1975 ? done_flag2 : c1976 ? done_flag2 : c1977 ? done_flag2 : c1978 ? done_flag2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? exec_result336 : (((c2019 || c2017) || c2018) || c2016) ? exec_result346 : c1981 ? done_flag2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? exec_result357 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? exec_result367 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? exec_result377 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? exec_result387 : (((c2038 || c2040) || c2037) || c2039) ? exec_result396 : (c2041 || c2042) ? exec_result404 : c1988 ? done_flag2 : c1989 ? done_flag2 : c1990 ? done_flag2 : c1991 ? done_flag2 : c1992 ? done_flag2 : c1993 ? done_flag2 : c1994 ? done_flag2 : c1995 ? done_flag2 : c1996 ? done_flag2 : ((c2055 || c2091) || c2090) ? exec_result545 : c1998 ? done_flag2 : c1999 ? done_flag2 : c2000 ? done_flag2 : c2001 ? done_flag2 : (c2199 || c2198) ? done_flag2 : (c2002 && !c927) ? done_flag2 : c1972 ? done_flag2 : 'bz; */
          /* ip16 <= (c1971 && c889) ? ip2 : ((c2004 || c2005) || c2006) ? lit0_ip4 : c1974 ? ip2 : c1975 ? ip2 : c1976 ? ip2 : c1977 ? ip2 : c1978 ? ip2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? loop0_ip5 : (((c2019 || c2017) || c2018) || c2016) ? jump0_ip5 : c1981 ? address0_top2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? jump_ge0_ip5 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? jump_le0_ip5 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? jump_ne0_ip5 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? jump_eq0_ip5 : (((c2038 || c2040) || c2037) || c2039) ? point0_ip5 : (c2041 || c2042) ? write_point0_ip4 : c1988 ? ip2 : c1989 ? ip2 : c1990 ? ip2 : c1991 ? ip2 : c1992 ? ip2 : c1993 ? ip2 : c1994 ? ip2 : c1995 ? ip2 : c1996 ? ip2 : ((c2055 || c2091) || c2090) ? zero_pop_return0_ip5 : c1998 ? ip2 : c1999 ? ip2 : c2000 ? ip2 : c2001 ? ip2 : (c2199 || c2198) ? ip_inl554 : (c2002 && !c927) ? ip2 : c1972 ? ip15 : 'bz; */
          /* jump0_ip6 <= (c1971 && c889) ? jump0_ip2 : ((c2004 || c2005) || c2006) ? jump0_ip2 : c1974 ? jump0_ip2 : c1975 ? jump0_ip2 : c1976 ? jump0_ip2 : c1977 ? jump0_ip2 : c1978 ? jump0_ip2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? jump0_ip2 : (((c2019 || c2017) || c2018) || c2016) ? jump0_ip5 : c1981 ? jump0_ip2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? jump0_ip2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? jump0_ip2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? jump0_ip2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? jump0_ip2 : (((c2038 || c2040) || c2037) || c2039) ? jump0_ip2 : (c2041 || c2042) ? jump0_ip2 : c1988 ? jump0_ip2 : c1989 ? jump0_ip2 : c1990 ? jump0_ip2 : c1991 ? jump0_ip2 : c1992 ? jump0_ip2 : c1993 ? jump0_ip2 : c1994 ? jump0_ip2 : c1995 ? jump0_ip2 : c1996 ? jump0_ip2 : ((c2055 || c2091) || c2090) ? jump0_ip2 : c1998 ? jump0_ip2 : c1999 ? jump0_ip2 : c2000 ? jump0_ip2 : c2001 ? jump0_ip2 : (c2199 || c2198) ? jump0_ip2 : (c2002 && !c927) ? jump0_ip2 : c1972 ? jump0_ip2 : 'bz; */
          /* jump0_phase8 <= (c1971 && c889) ? jump0_phase2 : ((c2004 || c2005) || c2006) ? jump0_phase2 : c1974 ? jump0_phase2 : c1975 ? jump0_phase2 : c1976 ? jump0_phase2 : c1977 ? jump0_phase2 : c1978 ? jump0_phase2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? jump0_phase2 : (((c2019 || c2017) || c2018) || c2016) ? jump0_phase7 : c1981 ? jump0_phase2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? jump0_phase2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? jump0_phase2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? jump0_phase2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? jump0_phase2 : (((c2038 || c2040) || c2037) || c2039) ? jump0_phase2 : (c2041 || c2042) ? jump0_phase2 : c1988 ? jump0_phase2 : c1989 ? jump0_phase2 : c1990 ? jump0_phase2 : c1991 ? jump0_phase2 : c1992 ? jump0_phase2 : c1993 ? jump0_phase2 : c1994 ? jump0_phase2 : c1995 ? jump0_phase2 : c1996 ? jump0_phase2 : ((c2055 || c2091) || c2090) ? jump0_phase2 : c1998 ? jump0_phase2 : c1999 ? jump0_phase2 : c2000 ? jump0_phase2 : c2001 ? jump0_phase2 : (c2199 || c2198) ? jump0_phase2 : (c2002 && !c927) ? jump0_phase2 : c1972 ? jump0_phase2 : 'bz; */
          /* jump_eq0_a5 <= (c1971 && c889) ? jump_eq0_a2 : ((c2004 || c2005) || c2006) ? jump_eq0_a2 : c1974 ? jump_eq0_a2 : c1975 ? jump_eq0_a2 : c1976 ? jump_eq0_a2 : c1977 ? jump_eq0_a2 : c1978 ? jump_eq0_a2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? jump_eq0_a2 : (((c2019 || c2017) || c2018) || c2016) ? jump_eq0_a2 : c1981 ? jump_eq0_a2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? jump_eq0_a2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? jump_eq0_a2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? jump_eq0_a2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? jump_eq0_a4 : (((c2038 || c2040) || c2037) || c2039) ? jump_eq0_a2 : (c2041 || c2042) ? jump_eq0_a2 : c1988 ? jump_eq0_a2 : c1989 ? jump_eq0_a2 : c1990 ? jump_eq0_a2 : c1991 ? jump_eq0_a2 : c1992 ? jump_eq0_a2 : c1993 ? jump_eq0_a2 : c1994 ? jump_eq0_a2 : c1995 ? jump_eq0_a2 : c1996 ? jump_eq0_a2 : ((c2055 || c2091) || c2090) ? jump_eq0_a2 : c1998 ? jump_eq0_a2 : c1999 ? jump_eq0_a2 : c2000 ? jump_eq0_a2 : c2001 ? jump_eq0_a2 : (c2199 || c2198) ? jump_eq0_a2 : (c2002 && !c927) ? jump_eq0_a2 : c1972 ? jump_eq0_a2 : 'bz; */
          /* jump_eq0_ip6 <= (c1971 && c889) ? jump_eq0_ip2 : ((c2004 || c2005) || c2006) ? jump_eq0_ip2 : c1974 ? jump_eq0_ip2 : c1975 ? jump_eq0_ip2 : c1976 ? jump_eq0_ip2 : c1977 ? jump_eq0_ip2 : c1978 ? jump_eq0_ip2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? jump_eq0_ip2 : (((c2019 || c2017) || c2018) || c2016) ? jump_eq0_ip2 : c1981 ? jump_eq0_ip2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? jump_eq0_ip2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? jump_eq0_ip2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? jump_eq0_ip2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? jump_eq0_ip5 : (((c2038 || c2040) || c2037) || c2039) ? jump_eq0_ip2 : (c2041 || c2042) ? jump_eq0_ip2 : c1988 ? jump_eq0_ip2 : c1989 ? jump_eq0_ip2 : c1990 ? jump_eq0_ip2 : c1991 ? jump_eq0_ip2 : c1992 ? jump_eq0_ip2 : c1993 ? jump_eq0_ip2 : c1994 ? jump_eq0_ip2 : c1995 ? jump_eq0_ip2 : c1996 ? jump_eq0_ip2 : ((c2055 || c2091) || c2090) ? jump_eq0_ip2 : c1998 ? jump_eq0_ip2 : c1999 ? jump_eq0_ip2 : c2000 ? jump_eq0_ip2 : c2001 ? jump_eq0_ip2 : (c2199 || c2198) ? jump_eq0_ip2 : (c2002 && !c927) ? jump_eq0_ip2 : c1972 ? jump_eq0_ip2 : 'bz; */
          /* jump_eq0_phase9 <= (c1971 && c889) ? jump_eq0_phase2 : ((c2004 || c2005) || c2006) ? jump_eq0_phase2 : c1974 ? jump_eq0_phase2 : c1975 ? jump_eq0_phase2 : c1976 ? jump_eq0_phase2 : c1977 ? jump_eq0_phase2 : c1978 ? jump_eq0_phase2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? jump_eq0_phase2 : (((c2019 || c2017) || c2018) || c2016) ? jump_eq0_phase2 : c1981 ? jump_eq0_phase2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? jump_eq0_phase2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? jump_eq0_phase2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? jump_eq0_phase2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? jump_eq0_phase8 : (((c2038 || c2040) || c2037) || c2039) ? jump_eq0_phase2 : (c2041 || c2042) ? jump_eq0_phase2 : c1988 ? jump_eq0_phase2 : c1989 ? jump_eq0_phase2 : c1990 ? jump_eq0_phase2 : c1991 ? jump_eq0_phase2 : c1992 ? jump_eq0_phase2 : c1993 ? jump_eq0_phase2 : c1994 ? jump_eq0_phase2 : c1995 ? jump_eq0_phase2 : c1996 ? jump_eq0_phase2 : ((c2055 || c2091) || c2090) ? jump_eq0_phase2 : c1998 ? jump_eq0_phase2 : c1999 ? jump_eq0_phase2 : c2000 ? jump_eq0_phase2 : c2001 ? jump_eq0_phase2 : (c2199 || c2198) ? jump_eq0_phase2 : (c2002 && !c927) ? jump_eq0_phase2 : c1972 ? jump_eq0_phase2 : 'bz; */
          /* jump_ge0_a5 <= (c1971 && c889) ? jump_ge0_a2 : ((c2004 || c2005) || c2006) ? jump_ge0_a2 : c1974 ? jump_ge0_a2 : c1975 ? jump_ge0_a2 : c1976 ? jump_ge0_a2 : c1977 ? jump_ge0_a2 : c1978 ? jump_ge0_a2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? jump_ge0_a2 : (((c2019 || c2017) || c2018) || c2016) ? jump_ge0_a2 : c1981 ? jump_ge0_a2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? jump_ge0_a4 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? jump_ge0_a2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? jump_ge0_a2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? jump_ge0_a2 : (((c2038 || c2040) || c2037) || c2039) ? jump_ge0_a2 : (c2041 || c2042) ? jump_ge0_a2 : c1988 ? jump_ge0_a2 : c1989 ? jump_ge0_a2 : c1990 ? jump_ge0_a2 : c1991 ? jump_ge0_a2 : c1992 ? jump_ge0_a2 : c1993 ? jump_ge0_a2 : c1994 ? jump_ge0_a2 : c1995 ? jump_ge0_a2 : c1996 ? jump_ge0_a2 : ((c2055 || c2091) || c2090) ? jump_ge0_a2 : c1998 ? jump_ge0_a2 : c1999 ? jump_ge0_a2 : c2000 ? jump_ge0_a2 : c2001 ? jump_ge0_a2 : (c2199 || c2198) ? jump_ge0_a2 : (c2002 && !c927) ? jump_ge0_a2 : c1972 ? jump_ge0_a2 : 'bz; */
          /* jump_ge0_ip6 <= (c1971 && c889) ? jump_ge0_ip2 : ((c2004 || c2005) || c2006) ? jump_ge0_ip2 : c1974 ? jump_ge0_ip2 : c1975 ? jump_ge0_ip2 : c1976 ? jump_ge0_ip2 : c1977 ? jump_ge0_ip2 : c1978 ? jump_ge0_ip2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? jump_ge0_ip2 : (((c2019 || c2017) || c2018) || c2016) ? jump_ge0_ip2 : c1981 ? jump_ge0_ip2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? jump_ge0_ip5 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? jump_ge0_ip2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? jump_ge0_ip2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? jump_ge0_ip2 : (((c2038 || c2040) || c2037) || c2039) ? jump_ge0_ip2 : (c2041 || c2042) ? jump_ge0_ip2 : c1988 ? jump_ge0_ip2 : c1989 ? jump_ge0_ip2 : c1990 ? jump_ge0_ip2 : c1991 ? jump_ge0_ip2 : c1992 ? jump_ge0_ip2 : c1993 ? jump_ge0_ip2 : c1994 ? jump_ge0_ip2 : c1995 ? jump_ge0_ip2 : c1996 ? jump_ge0_ip2 : ((c2055 || c2091) || c2090) ? jump_ge0_ip2 : c1998 ? jump_ge0_ip2 : c1999 ? jump_ge0_ip2 : c2000 ? jump_ge0_ip2 : c2001 ? jump_ge0_ip2 : (c2199 || c2198) ? jump_ge0_ip2 : (c2002 && !c927) ? jump_ge0_ip2 : c1972 ? jump_ge0_ip2 : 'bz; */
          /* jump_ge0_phase9 <= (c1971 && c889) ? jump_ge0_phase2 : ((c2004 || c2005) || c2006) ? jump_ge0_phase2 : c1974 ? jump_ge0_phase2 : c1975 ? jump_ge0_phase2 : c1976 ? jump_ge0_phase2 : c1977 ? jump_ge0_phase2 : c1978 ? jump_ge0_phase2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? jump_ge0_phase2 : (((c2019 || c2017) || c2018) || c2016) ? jump_ge0_phase2 : c1981 ? jump_ge0_phase2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? jump_ge0_phase8 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? jump_ge0_phase2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? jump_ge0_phase2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? jump_ge0_phase2 : (((c2038 || c2040) || c2037) || c2039) ? jump_ge0_phase2 : (c2041 || c2042) ? jump_ge0_phase2 : c1988 ? jump_ge0_phase2 : c1989 ? jump_ge0_phase2 : c1990 ? jump_ge0_phase2 : c1991 ? jump_ge0_phase2 : c1992 ? jump_ge0_phase2 : c1993 ? jump_ge0_phase2 : c1994 ? jump_ge0_phase2 : c1995 ? jump_ge0_phase2 : c1996 ? jump_ge0_phase2 : ((c2055 || c2091) || c2090) ? jump_ge0_phase2 : c1998 ? jump_ge0_phase2 : c1999 ? jump_ge0_phase2 : c2000 ? jump_ge0_phase2 : c2001 ? jump_ge0_phase2 : (c2199 || c2198) ? jump_ge0_phase2 : (c2002 && !c927) ? jump_ge0_phase2 : c1972 ? jump_ge0_phase2 : 'bz; */
          /* jump_le0_a5 <= (c1971 && c889) ? jump_le0_a2 : ((c2004 || c2005) || c2006) ? jump_le0_a2 : c1974 ? jump_le0_a2 : c1975 ? jump_le0_a2 : c1976 ? jump_le0_a2 : c1977 ? jump_le0_a2 : c1978 ? jump_le0_a2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? jump_le0_a2 : (((c2019 || c2017) || c2018) || c2016) ? jump_le0_a2 : c1981 ? jump_le0_a2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? jump_le0_a2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? jump_le0_a4 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? jump_le0_a2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? jump_le0_a2 : (((c2038 || c2040) || c2037) || c2039) ? jump_le0_a2 : (c2041 || c2042) ? jump_le0_a2 : c1988 ? jump_le0_a2 : c1989 ? jump_le0_a2 : c1990 ? jump_le0_a2 : c1991 ? jump_le0_a2 : c1992 ? jump_le0_a2 : c1993 ? jump_le0_a2 : c1994 ? jump_le0_a2 : c1995 ? jump_le0_a2 : c1996 ? jump_le0_a2 : ((c2055 || c2091) || c2090) ? jump_le0_a2 : c1998 ? jump_le0_a2 : c1999 ? jump_le0_a2 : c2000 ? jump_le0_a2 : c2001 ? jump_le0_a2 : (c2199 || c2198) ? jump_le0_a2 : (c2002 && !c927) ? jump_le0_a2 : c1972 ? jump_le0_a2 : 'bz; */
          /* jump_le0_ip6 <= (c1971 && c889) ? jump_le0_ip2 : ((c2004 || c2005) || c2006) ? jump_le0_ip2 : c1974 ? jump_le0_ip2 : c1975 ? jump_le0_ip2 : c1976 ? jump_le0_ip2 : c1977 ? jump_le0_ip2 : c1978 ? jump_le0_ip2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? jump_le0_ip2 : (((c2019 || c2017) || c2018) || c2016) ? jump_le0_ip2 : c1981 ? jump_le0_ip2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? jump_le0_ip2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? jump_le0_ip5 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? jump_le0_ip2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? jump_le0_ip2 : (((c2038 || c2040) || c2037) || c2039) ? jump_le0_ip2 : (c2041 || c2042) ? jump_le0_ip2 : c1988 ? jump_le0_ip2 : c1989 ? jump_le0_ip2 : c1990 ? jump_le0_ip2 : c1991 ? jump_le0_ip2 : c1992 ? jump_le0_ip2 : c1993 ? jump_le0_ip2 : c1994 ? jump_le0_ip2 : c1995 ? jump_le0_ip2 : c1996 ? jump_le0_ip2 : ((c2055 || c2091) || c2090) ? jump_le0_ip2 : c1998 ? jump_le0_ip2 : c1999 ? jump_le0_ip2 : c2000 ? jump_le0_ip2 : c2001 ? jump_le0_ip2 : (c2199 || c2198) ? jump_le0_ip2 : (c2002 && !c927) ? jump_le0_ip2 : c1972 ? jump_le0_ip2 : 'bz; */
          /* jump_le0_phase9 <= (c1971 && c889) ? jump_le0_phase2 : ((c2004 || c2005) || c2006) ? jump_le0_phase2 : c1974 ? jump_le0_phase2 : c1975 ? jump_le0_phase2 : c1976 ? jump_le0_phase2 : c1977 ? jump_le0_phase2 : c1978 ? jump_le0_phase2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? jump_le0_phase2 : (((c2019 || c2017) || c2018) || c2016) ? jump_le0_phase2 : c1981 ? jump_le0_phase2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? jump_le0_phase2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? jump_le0_phase8 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? jump_le0_phase2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? jump_le0_phase2 : (((c2038 || c2040) || c2037) || c2039) ? jump_le0_phase2 : (c2041 || c2042) ? jump_le0_phase2 : c1988 ? jump_le0_phase2 : c1989 ? jump_le0_phase2 : c1990 ? jump_le0_phase2 : c1991 ? jump_le0_phase2 : c1992 ? jump_le0_phase2 : c1993 ? jump_le0_phase2 : c1994 ? jump_le0_phase2 : c1995 ? jump_le0_phase2 : c1996 ? jump_le0_phase2 : ((c2055 || c2091) || c2090) ? jump_le0_phase2 : c1998 ? jump_le0_phase2 : c1999 ? jump_le0_phase2 : c2000 ? jump_le0_phase2 : c2001 ? jump_le0_phase2 : (c2199 || c2198) ? jump_le0_phase2 : (c2002 && !c927) ? jump_le0_phase2 : c1972 ? jump_le0_phase2 : 'bz; */
          /* jump_ne0_a5 <= (c1971 && c889) ? jump_ne0_a2 : ((c2004 || c2005) || c2006) ? jump_ne0_a2 : c1974 ? jump_ne0_a2 : c1975 ? jump_ne0_a2 : c1976 ? jump_ne0_a2 : c1977 ? jump_ne0_a2 : c1978 ? jump_ne0_a2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? jump_ne0_a2 : (((c2019 || c2017) || c2018) || c2016) ? jump_ne0_a2 : c1981 ? jump_ne0_a2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? jump_ne0_a2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? jump_ne0_a2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? jump_ne0_a4 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? jump_ne0_a2 : (((c2038 || c2040) || c2037) || c2039) ? jump_ne0_a2 : (c2041 || c2042) ? jump_ne0_a2 : c1988 ? jump_ne0_a2 : c1989 ? jump_ne0_a2 : c1990 ? jump_ne0_a2 : c1991 ? jump_ne0_a2 : c1992 ? jump_ne0_a2 : c1993 ? jump_ne0_a2 : c1994 ? jump_ne0_a2 : c1995 ? jump_ne0_a2 : c1996 ? jump_ne0_a2 : ((c2055 || c2091) || c2090) ? jump_ne0_a2 : c1998 ? jump_ne0_a2 : c1999 ? jump_ne0_a2 : c2000 ? jump_ne0_a2 : c2001 ? jump_ne0_a2 : (c2199 || c2198) ? jump_ne0_a2 : (c2002 && !c927) ? jump_ne0_a2 : c1972 ? jump_ne0_a2 : 'bz; */
          /* jump_ne0_ip6 <= (c1971 && c889) ? jump_ne0_ip2 : ((c2004 || c2005) || c2006) ? jump_ne0_ip2 : c1974 ? jump_ne0_ip2 : c1975 ? jump_ne0_ip2 : c1976 ? jump_ne0_ip2 : c1977 ? jump_ne0_ip2 : c1978 ? jump_ne0_ip2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? jump_ne0_ip2 : (((c2019 || c2017) || c2018) || c2016) ? jump_ne0_ip2 : c1981 ? jump_ne0_ip2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? jump_ne0_ip2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? jump_ne0_ip2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? jump_ne0_ip5 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? jump_ne0_ip2 : (((c2038 || c2040) || c2037) || c2039) ? jump_ne0_ip2 : (c2041 || c2042) ? jump_ne0_ip2 : c1988 ? jump_ne0_ip2 : c1989 ? jump_ne0_ip2 : c1990 ? jump_ne0_ip2 : c1991 ? jump_ne0_ip2 : c1992 ? jump_ne0_ip2 : c1993 ? jump_ne0_ip2 : c1994 ? jump_ne0_ip2 : c1995 ? jump_ne0_ip2 : c1996 ? jump_ne0_ip2 : ((c2055 || c2091) || c2090) ? jump_ne0_ip2 : c1998 ? jump_ne0_ip2 : c1999 ? jump_ne0_ip2 : c2000 ? jump_ne0_ip2 : c2001 ? jump_ne0_ip2 : (c2199 || c2198) ? jump_ne0_ip2 : (c2002 && !c927) ? jump_ne0_ip2 : c1972 ? jump_ne0_ip2 : 'bz; */
          /* jump_ne0_phase9 <= (c1971 && c889) ? jump_ne0_phase2 : ((c2004 || c2005) || c2006) ? jump_ne0_phase2 : c1974 ? jump_ne0_phase2 : c1975 ? jump_ne0_phase2 : c1976 ? jump_ne0_phase2 : c1977 ? jump_ne0_phase2 : c1978 ? jump_ne0_phase2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? jump_ne0_phase2 : (((c2019 || c2017) || c2018) || c2016) ? jump_ne0_phase2 : c1981 ? jump_ne0_phase2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? jump_ne0_phase2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? jump_ne0_phase2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? jump_ne0_phase8 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? jump_ne0_phase2 : (((c2038 || c2040) || c2037) || c2039) ? jump_ne0_phase2 : (c2041 || c2042) ? jump_ne0_phase2 : c1988 ? jump_ne0_phase2 : c1989 ? jump_ne0_phase2 : c1990 ? jump_ne0_phase2 : c1991 ? jump_ne0_phase2 : c1992 ? jump_ne0_phase2 : c1993 ? jump_ne0_phase2 : c1994 ? jump_ne0_phase2 : c1995 ? jump_ne0_phase2 : c1996 ? jump_ne0_phase2 : ((c2055 || c2091) || c2090) ? jump_ne0_phase2 : c1998 ? jump_ne0_phase2 : c1999 ? jump_ne0_phase2 : c2000 ? jump_ne0_phase2 : c2001 ? jump_ne0_phase2 : (c2199 || c2198) ? jump_ne0_phase2 : (c2002 && !c927) ? jump_ne0_phase2 : c1972 ? jump_ne0_phase2 : 'bz; */
          /* lit0_ip5 <= (c1971 && c889) ? lit0_ip2 : ((c2004 || c2005) || c2006) ? lit0_ip4 : c1974 ? lit0_ip2 : c1975 ? lit0_ip2 : c1976 ? lit0_ip2 : c1977 ? lit0_ip2 : c1978 ? lit0_ip2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? lit0_ip2 : (((c2019 || c2017) || c2018) || c2016) ? lit0_ip2 : c1981 ? lit0_ip2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? lit0_ip2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? lit0_ip2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? lit0_ip2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? lit0_ip2 : (((c2038 || c2040) || c2037) || c2039) ? lit0_ip2 : (c2041 || c2042) ? lit0_ip2 : c1988 ? lit0_ip2 : c1989 ? lit0_ip2 : c1990 ? lit0_ip2 : c1991 ? lit0_ip2 : c1992 ? lit0_ip2 : c1993 ? lit0_ip2 : c1994 ? lit0_ip2 : c1995 ? lit0_ip2 : c1996 ? lit0_ip2 : ((c2055 || c2091) || c2090) ? lit0_ip2 : c1998 ? lit0_ip2 : c1999 ? lit0_ip2 : c2000 ? lit0_ip2 : c2001 ? lit0_ip2 : (c2199 || c2198) ? lit0_ip2 : (c2002 && !c927) ? lit0_ip2 : c1972 ? lit0_ip2 : 'bz; */
          /* lit0_phase7 <= (c1971 && c889) ? lit0_phase2 : ((c2004 || c2005) || c2006) ? lit0_phase6 : c1974 ? lit0_phase2 : c1975 ? lit0_phase2 : c1976 ? lit0_phase2 : c1977 ? lit0_phase2 : c1978 ? lit0_phase2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? lit0_phase2 : (((c2019 || c2017) || c2018) || c2016) ? lit0_phase2 : c1981 ? lit0_phase2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? lit0_phase2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? lit0_phase2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? lit0_phase2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? lit0_phase2 : (((c2038 || c2040) || c2037) || c2039) ? lit0_phase2 : (c2041 || c2042) ? lit0_phase2 : c1988 ? lit0_phase2 : c1989 ? lit0_phase2 : c1990 ? lit0_phase2 : c1991 ? lit0_phase2 : c1992 ? lit0_phase2 : c1993 ? lit0_phase2 : c1994 ? lit0_phase2 : c1995 ? lit0_phase2 : c1996 ? lit0_phase2 : ((c2055 || c2091) || c2090) ? lit0_phase2 : c1998 ? lit0_phase2 : c1999 ? lit0_phase2 : c2000 ? lit0_phase2 : c2001 ? lit0_phase2 : (c2199 || c2198) ? lit0_phase2 : (c2002 && !c927) ? lit0_phase2 : c1972 ? lit0_phase2 : 'bz; */
          /* loop0_ip6 <= (c1971 && c889) ? loop0_ip2 : ((c2004 || c2005) || c2006) ? loop0_ip2 : c1974 ? loop0_ip2 : c1975 ? loop0_ip2 : c1976 ? loop0_ip2 : c1977 ? loop0_ip2 : c1978 ? loop0_ip2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? loop0_ip5 : (((c2019 || c2017) || c2018) || c2016) ? loop0_ip2 : c1981 ? loop0_ip2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? loop0_ip2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? loop0_ip2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? loop0_ip2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? loop0_ip2 : (((c2038 || c2040) || c2037) || c2039) ? loop0_ip2 : (c2041 || c2042) ? loop0_ip2 : c1988 ? loop0_ip2 : c1989 ? loop0_ip2 : c1990 ? loop0_ip2 : c1991 ? loop0_ip2 : c1992 ? loop0_ip2 : c1993 ? loop0_ip2 : c1994 ? loop0_ip2 : c1995 ? loop0_ip2 : c1996 ? loop0_ip2 : ((c2055 || c2091) || c2090) ? loop0_ip2 : c1998 ? loop0_ip2 : c1999 ? loop0_ip2 : c2000 ? loop0_ip2 : c2001 ? loop0_ip2 : (c2199 || c2198) ? loop0_ip2 : (c2002 && !c927) ? loop0_ip2 : c1972 ? loop0_ip2 : 'bz; */
          /* loop0_phase9 <= (c1971 && c889) ? loop0_phase2 : ((c2004 || c2005) || c2006) ? loop0_phase2 : c1974 ? loop0_phase2 : c1975 ? loop0_phase2 : c1976 ? loop0_phase2 : c1977 ? loop0_phase2 : c1978 ? loop0_phase2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? loop0_phase8 : (((c2019 || c2017) || c2018) || c2016) ? loop0_phase2 : c1981 ? loop0_phase2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? loop0_phase2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? loop0_phase2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? loop0_phase2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? loop0_phase2 : (((c2038 || c2040) || c2037) || c2039) ? loop0_phase2 : (c2041 || c2042) ? loop0_phase2 : c1988 ? loop0_phase2 : c1989 ? loop0_phase2 : c1990 ? loop0_phase2 : c1991 ? loop0_phase2 : c1992 ? loop0_phase2 : c1993 ? loop0_phase2 : c1994 ? loop0_phase2 : c1995 ? loop0_phase2 : c1996 ? loop0_phase2 : ((c2055 || c2091) || c2090) ? loop0_phase2 : c1998 ? loop0_phase2 : c1999 ? loop0_phase2 : c2000 ? loop0_phase2 : c2001 ? loop0_phase2 : (c2199 || c2198) ? loop0_phase2 : (c2002 && !c927) ? loop0_phase2 : c1972 ? loop0_phase2 : 'bz; */
          /* point0_ip6 <= (c1971 && c889) ? point0_ip2 : ((c2004 || c2005) || c2006) ? point0_ip2 : c1974 ? point0_ip2 : c1975 ? point0_ip2 : c1976 ? point0_ip2 : c1977 ? point0_ip2 : c1978 ? point0_ip2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? point0_ip2 : (((c2019 || c2017) || c2018) || c2016) ? point0_ip2 : c1981 ? point0_ip2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? point0_ip2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? point0_ip2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? point0_ip2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? point0_ip2 : (((c2038 || c2040) || c2037) || c2039) ? point0_ip5 : (c2041 || c2042) ? point0_ip2 : c1988 ? point0_ip2 : c1989 ? point0_ip2 : c1990 ? point0_ip2 : c1991 ? point0_ip2 : c1992 ? point0_ip2 : c1993 ? point0_ip2 : c1994 ? point0_ip2 : c1995 ? point0_ip2 : c1996 ? point0_ip2 : ((c2055 || c2091) || c2090) ? point0_ip2 : c1998 ? point0_ip2 : c1999 ? point0_ip2 : c2000 ? point0_ip2 : c2001 ? point0_ip2 : (c2199 || c2198) ? point0_ip2 : (c2002 && !c927) ? point0_ip2 : c1972 ? point0_ip2 : 'bz; */
          /* point0_ip_saved5 <= (c1971 && c889) ? point0_ip_saved2 : ((c2004 || c2005) || c2006) ? point0_ip_saved2 : c1974 ? point0_ip_saved2 : c1975 ? point0_ip_saved2 : c1976 ? point0_ip_saved2 : c1977 ? point0_ip_saved2 : c1978 ? point0_ip_saved2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? point0_ip_saved2 : (((c2019 || c2017) || c2018) || c2016) ? point0_ip_saved2 : c1981 ? point0_ip_saved2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? point0_ip_saved2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? point0_ip_saved2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? point0_ip_saved2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? point0_ip_saved2 : (((c2038 || c2040) || c2037) || c2039) ? point0_ip_saved4 : (c2041 || c2042) ? point0_ip_saved2 : c1988 ? point0_ip_saved2 : c1989 ? point0_ip_saved2 : c1990 ? point0_ip_saved2 : c1991 ? point0_ip_saved2 : c1992 ? point0_ip_saved2 : c1993 ? point0_ip_saved2 : c1994 ? point0_ip_saved2 : c1995 ? point0_ip_saved2 : c1996 ? point0_ip_saved2 : ((c2055 || c2091) || c2090) ? point0_ip_saved2 : c1998 ? point0_ip_saved2 : c1999 ? point0_ip_saved2 : c2000 ? point0_ip_saved2 : c2001 ? point0_ip_saved2 : (c2199 || c2198) ? point0_ip_saved2 : (c2002 && !c927) ? point0_ip_saved2 : c1972 ? point0_ip_saved2 : 'bz; */
          /* point0_phase8 <= (c1971 && c889) ? point0_phase2 : ((c2004 || c2005) || c2006) ? point0_phase2 : c1974 ? point0_phase2 : c1975 ? point0_phase2 : c1976 ? point0_phase2 : c1977 ? point0_phase2 : c1978 ? point0_phase2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? point0_phase2 : (((c2019 || c2017) || c2018) || c2016) ? point0_phase2 : c1981 ? point0_phase2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? point0_phase2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? point0_phase2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? point0_phase2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? point0_phase2 : (((c2038 || c2040) || c2037) || c2039) ? point0_phase7 : (c2041 || c2042) ? point0_phase2 : c1988 ? point0_phase2 : c1989 ? point0_phase2 : c1990 ? point0_phase2 : c1991 ? point0_phase2 : c1992 ? point0_phase2 : c1993 ? point0_phase2 : c1994 ? point0_phase2 : c1995 ? point0_phase2 : c1996 ? point0_phase2 : ((c2055 || c2091) || c2090) ? point0_phase2 : c1998 ? point0_phase2 : c1999 ? point0_phase2 : c2000 ? point0_phase2 : c2001 ? point0_phase2 : (c2199 || c2198) ? point0_phase2 : (c2002 && !c927) ? point0_phase2 : c1972 ? point0_phase2 : 'bz; */
          /* stack0_pos43 <= (c1971 && c889) ? stack0_pos2 : ((c2004 || c2005) || c2006) ? stack0_pos4 : c1974 ? stack0_pos5 : c1975 ? stack0_pos6 : c1976 ? stack0_pos2 : c1977 ? stack0_pos7 : c1978 ? stack0_pos8 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? stack0_pos10 : (((c2019 || c2017) || c2018) || c2016) ? stack0_pos2 : c1981 ? stack0_pos2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? stack0_pos13 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? stack0_pos16 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? stack0_pos19 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? stack0_pos22 : (((c2038 || c2040) || c2037) || c2039) ? stack0_pos2 : (c2041 || c2042) ? stack0_pos25 : c1988 ? stack0_pos26 : c1989 ? stack0_pos27 : c1990 ? stack0_pos28 : c1991 ? stack0_pos2 : c1992 ? stack0_pos29 : c1993 ? stack0_pos30 : c1994 ? stack0_pos31 : c1995 ? stack0_pos32 : c1996 ? stack0_pos33 : ((c2055 || c2091) || c2090) ? stack0_pos35 : c1998 ? stack0_pos2 : c1999 ? stack0_pos2 : c2000 ? stack0_pos2 : c2001 ? stack0_pos37 : (c2199 || c2198) ? stack0_pos42 : (c2002 && !c927) ? stack0_pos2 : c1972 ? stack0_pos2 : 'bz; */
          /* stack0_second45 <= (c1971 && c889) ? stack0_second2 : ((c2004 || c2005) || c2006) ? stack0_second4 : c1974 ? stack0_top2 : c1975 ? stack0_second6 : c1976 ? stack0_top2 : c1977 ? stack0_second8 : c1978 ? stack0_top2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? stack0_second11 : (((c2019 || c2017) || c2018) || c2016) ? stack0_second2 : c1981 ? stack0_second2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? stack0_second14 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? stack0_second17 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? stack0_second20 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? stack0_second23 : (((c2038 || c2040) || c2037) || c2039) ? stack0_second2 : (c2041 || c2042) ? stack0_second26 : c1988 ? stack0_second27 : c1989 ? stack0_second28 : c1990 ? stack0_second29 : c1991 ? stack0_second30 : c1992 ? stack0_second31 : c1993 ? stack0_second32 : c1994 ? stack0_second33 : c1995 ? stack0_second34 : c1996 ? stack0_second35 : ((c2055 || c2091) || c2090) ? stack0_second37 : c1998 ? stack0_second2 : c1999 ? stack0_second2 : c2000 ? stack0_second2 : c2001 ? stack0_second39 : (c2199 || c2198) ? stack0_second44 : (c2002 && !c927) ? stack0_second2 : c1972 ? stack0_second2 : 'bz; */
          /* stack0_top59 <= (c1971 && c889) ? stack0_top2 : ((c2004 || c2005) || c2006) ? stack0_top4 : c1974 ? stack0_top2 : c1975 ? stack0_second2 : c1976 ? stack0_second2 : c1977 ? stack0_second2 : c1978 ? address0_top2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? stack0_top12 : (((c2019 || c2017) || c2018) || c2016) ? stack0_top2 : c1981 ? stack0_top2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? stack0_top15 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? stack0_top18 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? stack0_top21 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? stack0_top24 : (((c2038 || c2040) || c2037) || c2039) ? stack0_top26 : (c2041 || c2042) ? stack0_second2 : c1988 ? stack0_top31 : c1989 ? stack0_top33 : c1990 ? stack0_top35 : c1991 ? stack0_top36 : c1992 ? stack0_top38 : c1993 ? stack0_top40 : c1994 ? stack0_top42 : c1995 ? stack0_top44 : c1996 ? stack0_top46 : ((c2055 || c2091) || c2090) ? stack0_top48 : c1998 ? stack0_top49 : c1999 ? stack0_top50 : c2000 ? stack0_top51 : c2001 ? stack0_second38 : (c2199 || c2198) ? stack0_top58 : (c2002 && !c927) ? stack0_top2 : c1972 ? stack0_top2 : 'bz; */
          t11 <= (c1971 && c889) ? t11 : ((c2004 || c2005) || c2006) ? t11 : c1974 ? t11 : c1975 ? t11 : c1976 ? t11 : c1977 ? t11 : c1978 ? t11 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? t11 : (((c2019 || c2017) || c2018) || c2016) ? t11 : c1981 ? t11 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? t11 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? t11 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? t11 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? t11 : (((c2038 || c2040) || c2037) || c2039) ? t11 : (c2041 || c2042) ? t11 : c1988 ? stack0_top2 : c1989 ? stack0_top2 : c1990 ? stack0_top2 : c1991 ? t11 : c1992 ? stack0_top2 : c1993 ? stack0_top2 : c1994 ? stack0_top2 : c1995 ? stack0_top2 : c1996 ? stack0_top2 : ((c2055 || c2091) || c2090) ? t11 : c1998 ? t11 : c1999 ? t11 : c2000 ? stack0_top2 : c2001 ? t11 : (c2199 || c2198) ? t11 : (c2002 && !c927) ? t11 : c1972 ? t11 : 'bz;
          /* wr_flag4 <= (c1971 && c889) ? wr_flag2 : ((c2004 || c2005) || c2006) ? wr_flag2 : c1974 ? wr_flag2 : c1975 ? wr_flag2 : c1976 ? wr_flag2 : c1977 ? wr_flag2 : c1978 ? wr_flag2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? wr_flag2 : (((c2019 || c2017) || c2018) || c2016) ? wr_flag2 : c1981 ? wr_flag2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? wr_flag2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? wr_flag2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? wr_flag2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? wr_flag2 : (((c2038 || c2040) || c2037) || c2039) ? wr_flag2 : (c2041 || c2042) ? t2829 : c1988 ? wr_flag2 : c1989 ? wr_flag2 : c1990 ? wr_flag2 : c1991 ? wr_flag2 : c1992 ? wr_flag2 : c1993 ? wr_flag2 : c1994 ? wr_flag2 : c1995 ? wr_flag2 : c1996 ? wr_flag2 : ((c2055 || c2091) || c2090) ? wr_flag2 : c1998 ? wr_flag2 : c1999 ? wr_flag2 : c2000 ? wr_flag2 : c2001 ? wr_flag2 : (c2199 || c2198) ? wr_flag2 : (c2002 && !c927) ? wr_flag2 : c1972 ? wr_flag2 : 'bz; */
          /* wr_mem_addr4 <= (c1971 && c889) ? wr_mem_addr2 : ((c2004 || c2005) || c2006) ? wr_mem_addr2 : c1974 ? wr_mem_addr2 : c1975 ? wr_mem_addr2 : c1976 ? wr_mem_addr2 : c1977 ? wr_mem_addr2 : c1978 ? wr_mem_addr2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? wr_mem_addr2 : (((c2019 || c2017) || c2018) || c2016) ? wr_mem_addr2 : c1981 ? wr_mem_addr2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? wr_mem_addr2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? wr_mem_addr2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? wr_mem_addr2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? wr_mem_addr2 : (((c2038 || c2040) || c2037) || c2039) ? wr_mem_addr2 : (c2041 || c2042) ? t2830 : c1988 ? wr_mem_addr2 : c1989 ? wr_mem_addr2 : c1990 ? wr_mem_addr2 : c1991 ? wr_mem_addr2 : c1992 ? wr_mem_addr2 : c1993 ? wr_mem_addr2 : c1994 ? wr_mem_addr2 : c1995 ? wr_mem_addr2 : c1996 ? wr_mem_addr2 : ((c2055 || c2091) || c2090) ? wr_mem_addr2 : c1998 ? wr_mem_addr2 : c1999 ? wr_mem_addr2 : c2000 ? wr_mem_addr2 : c2001 ? wr_mem_addr2 : (c2199 || c2198) ? wr_mem_addr2 : (c2002 && !c927) ? wr_mem_addr2 : c1972 ? wr_mem_addr2 : 'bz; */
          /* wr_mem_data4 <= (c1971 && c889) ? wr_mem_data2 : ((c2004 || c2005) || c2006) ? wr_mem_data2 : c1974 ? wr_mem_data2 : c1975 ? wr_mem_data2 : c1976 ? wr_mem_data2 : c1977 ? wr_mem_data2 : c1978 ? wr_mem_data2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? wr_mem_data2 : (((c2019 || c2017) || c2018) || c2016) ? wr_mem_data2 : c1981 ? wr_mem_data2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? wr_mem_data2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? wr_mem_data2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? wr_mem_data2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? wr_mem_data2 : (((c2038 || c2040) || c2037) || c2039) ? wr_mem_data2 : (c2041 || c2042) ? t2831 : c1988 ? wr_mem_data2 : c1989 ? wr_mem_data2 : c1990 ? wr_mem_data2 : c1991 ? wr_mem_data2 : c1992 ? wr_mem_data2 : c1993 ? wr_mem_data2 : c1994 ? wr_mem_data2 : c1995 ? wr_mem_data2 : c1996 ? wr_mem_data2 : ((c2055 || c2091) || c2090) ? wr_mem_data2 : c1998 ? wr_mem_data2 : c1999 ? wr_mem_data2 : c2000 ? wr_mem_data2 : c2001 ? wr_mem_data2 : (c2199 || c2198) ? wr_mem_data2 : (c2002 && !c927) ? wr_mem_data2 : c1972 ? wr_mem_data2 : 'bz; */
          /* write_point0_addr5 <= (c1971 && c889) ? write_point0_addr2 : ((c2004 || c2005) || c2006) ? write_point0_addr2 : c1974 ? write_point0_addr2 : c1975 ? write_point0_addr2 : c1976 ? write_point0_addr2 : c1977 ? write_point0_addr2 : c1978 ? write_point0_addr2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? write_point0_addr2 : (((c2019 || c2017) || c2018) || c2016) ? write_point0_addr2 : c1981 ? write_point0_addr2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? write_point0_addr2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? write_point0_addr2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? write_point0_addr2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? write_point0_addr2 : (((c2038 || c2040) || c2037) || c2039) ? write_point0_addr2 : (c2041 || c2042) ? write_point0_addr4 : c1988 ? write_point0_addr2 : c1989 ? write_point0_addr2 : c1990 ? write_point0_addr2 : c1991 ? write_point0_addr2 : c1992 ? write_point0_addr2 : c1993 ? write_point0_addr2 : c1994 ? write_point0_addr2 : c1995 ? write_point0_addr2 : c1996 ? write_point0_addr2 : ((c2055 || c2091) || c2090) ? write_point0_addr2 : c1998 ? write_point0_addr2 : c1999 ? write_point0_addr2 : c2000 ? write_point0_addr2 : c2001 ? write_point0_addr2 : (c2199 || c2198) ? write_point0_addr2 : (c2002 && !c927) ? write_point0_addr2 : c1972 ? write_point0_addr2 : 'bz; */
          /* write_point0_data5 <= (c1971 && c889) ? write_point0_data2 : ((c2004 || c2005) || c2006) ? write_point0_data2 : c1974 ? write_point0_data2 : c1975 ? write_point0_data2 : c1976 ? write_point0_data2 : c1977 ? write_point0_data2 : c1978 ? write_point0_data2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? write_point0_data2 : (((c2019 || c2017) || c2018) || c2016) ? write_point0_data2 : c1981 ? write_point0_data2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? write_point0_data2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? write_point0_data2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? write_point0_data2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? write_point0_data2 : (((c2038 || c2040) || c2037) || c2039) ? write_point0_data2 : (c2041 || c2042) ? write_point0_data4 : c1988 ? write_point0_data2 : c1989 ? write_point0_data2 : c1990 ? write_point0_data2 : c1991 ? write_point0_data2 : c1992 ? write_point0_data2 : c1993 ? write_point0_data2 : c1994 ? write_point0_data2 : c1995 ? write_point0_data2 : c1996 ? write_point0_data2 : ((c2055 || c2091) || c2090) ? write_point0_data2 : c1998 ? write_point0_data2 : c1999 ? write_point0_data2 : c2000 ? write_point0_data2 : c2001 ? write_point0_data2 : (c2199 || c2198) ? write_point0_data2 : (c2002 && !c927) ? write_point0_data2 : c1972 ? write_point0_data2 : 'bz; */
          /* write_point0_ip5 <= (c1971 && c889) ? write_point0_ip2 : ((c2004 || c2005) || c2006) ? write_point0_ip2 : c1974 ? write_point0_ip2 : c1975 ? write_point0_ip2 : c1976 ? write_point0_ip2 : c1977 ? write_point0_ip2 : c1978 ? write_point0_ip2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? write_point0_ip2 : (((c2019 || c2017) || c2018) || c2016) ? write_point0_ip2 : c1981 ? write_point0_ip2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? write_point0_ip2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? write_point0_ip2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? write_point0_ip2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? write_point0_ip2 : (((c2038 || c2040) || c2037) || c2039) ? write_point0_ip2 : (c2041 || c2042) ? write_point0_ip4 : c1988 ? write_point0_ip2 : c1989 ? write_point0_ip2 : c1990 ? write_point0_ip2 : c1991 ? write_point0_ip2 : c1992 ? write_point0_ip2 : c1993 ? write_point0_ip2 : c1994 ? write_point0_ip2 : c1995 ? write_point0_ip2 : c1996 ? write_point0_ip2 : ((c2055 || c2091) || c2090) ? write_point0_ip2 : c1998 ? write_point0_ip2 : c1999 ? write_point0_ip2 : c2000 ? write_point0_ip2 : c2001 ? write_point0_ip2 : (c2199 || c2198) ? write_point0_ip2 : (c2002 && !c927) ? write_point0_ip2 : c1972 ? write_point0_ip2 : 'bz; */
          /* write_point0_phase6 <= (c1971 && c889) ? write_point0_phase2 : ((c2004 || c2005) || c2006) ? write_point0_phase2 : c1974 ? write_point0_phase2 : c1975 ? write_point0_phase2 : c1976 ? write_point0_phase2 : c1977 ? write_point0_phase2 : c1978 ? write_point0_phase2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? write_point0_phase2 : (((c2019 || c2017) || c2018) || c2016) ? write_point0_phase2 : c1981 ? write_point0_phase2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? write_point0_phase2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? write_point0_phase2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? write_point0_phase2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? write_point0_phase2 : (((c2038 || c2040) || c2037) || c2039) ? write_point0_phase2 : (c2041 || c2042) ? write_point0_phase5 : c1988 ? write_point0_phase2 : c1989 ? write_point0_phase2 : c1990 ? write_point0_phase2 : c1991 ? write_point0_phase2 : c1992 ? write_point0_phase2 : c1993 ? write_point0_phase2 : c1994 ? write_point0_phase2 : c1995 ? write_point0_phase2 : c1996 ? write_point0_phase2 : ((c2055 || c2091) || c2090) ? write_point0_phase2 : c1998 ? write_point0_phase2 : c1999 ? write_point0_phase2 : c2000 ? write_point0_phase2 : c2001 ? write_point0_phase2 : (c2199 || c2198) ? write_point0_phase2 : (c2002 && !c927) ? write_point0_phase2 : c1972 ? write_point0_phase2 : 'bz; */
          /* zero_pop_return0_ip6 <= (c1971 && c889) ? zero_pop_return0_ip2 : ((c2004 || c2005) || c2006) ? zero_pop_return0_ip2 : c1974 ? zero_pop_return0_ip2 : c1975 ? zero_pop_return0_ip2 : c1976 ? zero_pop_return0_ip2 : c1977 ? zero_pop_return0_ip2 : c1978 ? zero_pop_return0_ip2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? zero_pop_return0_ip2 : (((c2019 || c2017) || c2018) || c2016) ? zero_pop_return0_ip2 : c1981 ? zero_pop_return0_ip2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? zero_pop_return0_ip2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? zero_pop_return0_ip2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? zero_pop_return0_ip2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? zero_pop_return0_ip2 : (((c2038 || c2040) || c2037) || c2039) ? zero_pop_return0_ip2 : (c2041 || c2042) ? zero_pop_return0_ip2 : c1988 ? zero_pop_return0_ip2 : c1989 ? zero_pop_return0_ip2 : c1990 ? zero_pop_return0_ip2 : c1991 ? zero_pop_return0_ip2 : c1992 ? zero_pop_return0_ip2 : c1993 ? zero_pop_return0_ip2 : c1994 ? zero_pop_return0_ip2 : c1995 ? zero_pop_return0_ip2 : c1996 ? zero_pop_return0_ip2 : ((c2055 || c2091) || c2090) ? zero_pop_return0_ip5 : c1998 ? zero_pop_return0_ip2 : c1999 ? zero_pop_return0_ip2 : c2000 ? zero_pop_return0_ip2 : c2001 ? zero_pop_return0_ip2 : (c2199 || c2198) ? zero_pop_return0_ip2 : (c2002 && !c927) ? zero_pop_return0_ip2 : c1972 ? zero_pop_return0_ip2 : 'bz; */
          /* zero_pop_return0_phase6 <= (c1971 && c889) ? zero_pop_return0_phase2 : ((c2004 || c2005) || c2006) ? zero_pop_return0_phase2 : c1974 ? zero_pop_return0_phase2 : c1975 ? zero_pop_return0_phase2 : c1976 ? zero_pop_return0_phase2 : c1977 ? zero_pop_return0_phase2 : c1978 ? zero_pop_return0_phase2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? zero_pop_return0_phase2 : (((c2019 || c2017) || c2018) || c2016) ? zero_pop_return0_phase2 : c1981 ? zero_pop_return0_phase2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? zero_pop_return0_phase2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? zero_pop_return0_phase2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? zero_pop_return0_phase2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? zero_pop_return0_phase2 : (((c2038 || c2040) || c2037) || c2039) ? zero_pop_return0_phase2 : (c2041 || c2042) ? zero_pop_return0_phase2 : c1988 ? zero_pop_return0_phase2 : c1989 ? zero_pop_return0_phase2 : c1990 ? zero_pop_return0_phase2 : c1991 ? zero_pop_return0_phase2 : c1992 ? zero_pop_return0_phase2 : c1993 ? zero_pop_return0_phase2 : c1994 ? zero_pop_return0_phase2 : c1995 ? zero_pop_return0_phase2 : c1996 ? zero_pop_return0_phase2 : ((c2055 || c2091) || c2090) ? zero_pop_return0_phase5 : c1998 ? zero_pop_return0_phase2 : c1999 ? zero_pop_return0_phase2 : c2000 ? zero_pop_return0_phase2 : c2001 ? zero_pop_return0_phase2 : (c2199 || c2198) ? zero_pop_return0_phase2 : (c2002 && !c927) ? zero_pop_return0_phase2 : c1972 ? zero_pop_return0_phase2 : 'bz; */
          /* c920 <= (wr_flag4 != 0); */
          /* c2200 <= (c886 && c920); */
          retro_main_state <= retro_main_L1_b178_S1;
        end
      end
      retro_main_L1_ifelse221_S3: begin
        _stack_addr <= t839_inl1_inl13;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= stack0_second2;
        /* t839_inl1_inl13 <= (stack0_pos2 - 2); */
        retro_main_state <= retro_main_L1_ifelse221_S4;
      end
      retro_main_L1_ifelse221_S4: begin
        _stack_req <= 0;
        retro_main_state <= retro_main_L1_exit219_S0;
      end
      retro_main_L1_ifthen304_S3: begin
        /* stack0_top10 <= (stack0_top2 - 1); */
        /* c875_inl33 <= (stack0_top10 != 0); */
        /* c876_inl33 <= (stack0_top10 > -1); */
        /* c877_inl33 <= (c875_inl33 && c876_inl33); */
        if (c877_inl33) begin
          /* c3402 <= (c3372 && c877_inl33); */
          /* c2124 <= (c2012 && c877_inl33); */
          retro_main_state <= retro_main_L1_exit310_S0;
        end else begin
          /* c3403 <= (c3372 && !c877_inl33); */
          /* c2125 <= (c2012 && !c877_inl33); */
          retro_main_state <= retro_main_L1_ifelse311_S5;
        end
      end
      retro_main_L1_ifthen317_S7: begin
        /* loop0_ip4 <= (mem_data - 1); */
        retro_main_state <= retro_main_L1_exit310_S0;
      end
      retro_main_L1_ifthen328_S1: begin
        /* jump_ge0_ip3 <= (ip2 + 1); */
        retro_main_state <= retro_main_L1_ifthen328_S3;
      end
      retro_main_L1_ifthen328_S3: begin
        _stack_addr <= t842_inl1_inl35;
        _stack_we <= 0;
        _stack_req <= 1;
        /* stack0_pos11 <= (stack0_pos2 - 1); */
        /* t842_inl1_inl35 <= (stack0_pos11 - 2); */
        retro_main_state <= retro_main_L1_ifthen328_S4;
      end
      retro_main_L1_ifthen328_S4: begin
        /*wait for output of _stack*/
        retro_main_state <= retro_main_L1_ifthen328_S5;
      end
      retro_main_L1_ifthen328_S5: begin
        stack0_second12 <= _stack_q;
        _stack_req <= 0;
        retro_main_state <= retro_main_L1_exit333_S0;
      end
      retro_main_L1_ifthen334_S4: begin
        _stack_addr <= t842_inl2_inl35;
        _stack_we <= 0;
        _stack_req <= 1;
        /* stack0_pos12 <= (stack0_pos2 - 1); */
        /* t842_inl2_inl35 <= (stack0_pos12 - 2); */
        retro_main_state <= retro_main_L1_ifthen334_S5;
      end
      retro_main_L1_ifthen334_S5: begin
        /*wait for output of _stack*/
        retro_main_state <= retro_main_L1_ifthen334_S6;
      end
      retro_main_L1_ifthen334_S6: begin
        stack0_second13 <= _stack_q;
        _stack_req <= 0;
        retro_main_state <= retro_main_L1_b564_S0;
      end
      retro_main_L1_ifthen341_S7: begin
        /* jump_ge0_ip4 <= (mem_data - 1); */
        retro_main_state <= retro_main_L1_exit333_S0;
      end
      retro_main_L1_ifthen345_S1: begin
        /* jump_le0_ip3 <= (ip2 + 1); */
        retro_main_state <= retro_main_L1_ifthen345_S4;
      end
      retro_main_L1_ifthen345_S4: begin
        _stack_addr <= t842_inl1_inl36;
        _stack_we <= 0;
        _stack_req <= 1;
        /* stack0_pos14 <= (stack0_pos2 - 1); */
        /* t842_inl1_inl36 <= (stack0_pos14 - 2); */
        retro_main_state <= retro_main_L1_ifthen345_S5;
      end
      retro_main_L1_ifthen345_S5: begin
        /*wait for output of _stack*/
        retro_main_state <= retro_main_L1_ifthen345_S6;
      end
      retro_main_L1_ifthen345_S6: begin
        stack0_second15 <= _stack_q;
        _stack_req <= 0;
        retro_main_state <= retro_main_L1_exit350_S0;
      end
      retro_main_L1_ifthen351_S4: begin
        _stack_addr <= t842_inl2_inl36;
        _stack_we <= 0;
        _stack_req <= 1;
        /* stack0_pos15 <= (stack0_pos2 - 1); */
        /* t842_inl2_inl36 <= (stack0_pos15 - 2); */
        retro_main_state <= retro_main_L1_ifthen351_S5;
      end
      retro_main_L1_ifthen351_S5: begin
        /*wait for output of _stack*/
        retro_main_state <= retro_main_L1_ifthen351_S6;
      end
      retro_main_L1_ifthen351_S6: begin
        stack0_second16 <= _stack_q;
        _stack_req <= 0;
        retro_main_state <= retro_main_L1_b565_S0;
      end
      retro_main_L1_ifthen358_S7: begin
        /* jump_le0_ip4 <= (mem_data - 1); */
        retro_main_state <= retro_main_L1_exit350_S0;
      end
      retro_main_L1_ifthen362_S1: begin
        /* jump_ne0_ip3 <= (ip2 + 1); */
        retro_main_state <= retro_main_L1_ifthen362_S4;
      end
      retro_main_L1_ifthen362_S4: begin
        _stack_addr <= t842_inl1_inl37;
        _stack_we <= 0;
        _stack_req <= 1;
        /* stack0_pos17 <= (stack0_pos2 - 1); */
        /* t842_inl1_inl37 <= (stack0_pos17 - 2); */
        retro_main_state <= retro_main_L1_ifthen362_S5;
      end
      retro_main_L1_ifthen362_S5: begin
        /*wait for output of _stack*/
        retro_main_state <= retro_main_L1_ifthen362_S6;
      end
      retro_main_L1_ifthen362_S6: begin
        stack0_second18 <= _stack_q;
        _stack_req <= 0;
        retro_main_state <= retro_main_L1_exit367_S0;
      end
      retro_main_L1_ifthen368_S4: begin
        _stack_addr <= t842_inl2_inl37;
        _stack_we <= 0;
        _stack_req <= 1;
        /* stack0_pos18 <= (stack0_pos2 - 1); */
        /* t842_inl2_inl37 <= (stack0_pos18 - 2); */
        retro_main_state <= retro_main_L1_ifthen368_S5;
      end
      retro_main_L1_ifthen368_S5: begin
        /*wait for output of _stack*/
        retro_main_state <= retro_main_L1_ifthen368_S6;
      end
      retro_main_L1_ifthen368_S6: begin
        stack0_second19 <= _stack_q;
        _stack_req <= 0;
        retro_main_state <= retro_main_L1_b566_S0;
      end
      retro_main_L1_ifthen375_S7: begin
        /* jump_ne0_ip4 <= (mem_data - 1); */
        retro_main_state <= retro_main_L1_exit367_S0;
      end
      retro_main_L1_ifthen379_S1: begin
        /* jump_eq0_ip3 <= (ip2 + 1); */
        retro_main_state <= retro_main_L1_ifthen379_S5;
      end
      retro_main_L1_ifthen379_S5: begin
        _stack_addr <= t842_inl1_inl38;
        _stack_we <= 0;
        _stack_req <= 1;
        /* stack0_pos20 <= (stack0_pos2 - 1); */
        /* t842_inl1_inl38 <= (stack0_pos20 - 2); */
        retro_main_state <= retro_main_L1_ifthen379_S6;
      end
      retro_main_L1_ifthen379_S6: begin
        /*wait for output of _stack*/
        retro_main_state <= retro_main_L1_ifthen379_S7;
      end
      retro_main_L1_ifthen379_S7: begin
        stack0_second21 <= _stack_q;
        _stack_req <= 0;
        retro_main_state <= retro_main_L1_exit384_S0;
      end
      retro_main_L1_ifthen385_S5: begin
        _stack_addr <= t842_inl2_inl38;
        _stack_we <= 0;
        _stack_req <= 1;
        /* stack0_pos21 <= (stack0_pos2 - 1); */
        /* t842_inl2_inl38 <= (stack0_pos21 - 2); */
        retro_main_state <= retro_main_L1_ifthen385_S6;
      end
      retro_main_L1_ifthen385_S6: begin
        /*wait for output of _stack*/
        retro_main_state <= retro_main_L1_ifthen385_S7;
      end
      retro_main_L1_ifthen385_S7: begin
        stack0_second22 <= _stack_q;
        _stack_req <= 0;
        retro_main_state <= retro_main_L1_b567_S0;
      end
      retro_main_L1_ifthen392_S7: begin
        /* jump_eq0_ip4 <= (mem_data - 1); */
        retro_main_state <= retro_main_L1_exit384_S0;
      end
      retro_main_L1_ifthen407_S5: begin
        _stack_addr <= t842_inl1_inl40;
        _stack_we <= 0;
        _stack_req <= 1;
        /* stack0_pos23 <= (stack0_pos2 - 1); */
        /* t842_inl1_inl40 <= (stack0_pos23 - 2); */
        retro_main_state <= retro_main_L1_ifthen407_S6;
      end
      retro_main_L1_ifthen407_S6: begin
        /*wait for output of _stack*/
        retro_main_state <= retro_main_L1_ifthen407_S7;
      end
      retro_main_L1_ifthen407_S7: begin
        stack0_second24 <= _stack_q;
        _stack_req <= 0;
        retro_main_state <= retro_main_L1_exit412_S0;
      end
      retro_main_L1_ifelse413_S5: begin
        _stack_addr <= t842_inl2_inl40;
        _stack_we <= 0;
        _stack_req <= 1;
        /* stack0_pos24 <= (stack0_pos2 - 1); */
        /* t842_inl2_inl40 <= (stack0_pos24 - 2); */
        retro_main_state <= retro_main_L1_ifelse413_S6;
      end
      retro_main_L1_ifelse413_S6: begin
        /*wait for output of _stack*/
        retro_main_state <= retro_main_L1_ifelse413_S7;
      end
      retro_main_L1_ifelse413_S7: begin
        stack0_second25 <= _stack_q;
        _stack_req <= 0;
        retro_main_state <= retro_main_L1_exit412_S0;
      end
      retro_main_L1_ifthen140_S1: begin
        /* c930_inl55 <= (t929_inl55 == 1); */
        if (c930_inl55) begin
          /* c3407 <= (c3401 && c930_inl55); */
          /* c2093 <= (c2060 && c930_inl55); */
          $display("%s", "rx_chflush");
          $finish();
          retro_main_state <= retro_main_L1_ifthen493_S1;
        end else begin
          t934_inl55 <= array1010[2];
          /* c3409 <= (c3401 && !c930_inl55); */
          /* c2139 <= (c2060 && !c930_inl55); */
          /* c3410 <= (c3407 && !c933_inl55); */
          /* c2140 <= (c2093 && !c933_inl55); */
          retro_main_state <= retro_main_L1_b497_S1;
        end
      end
      retro_main_L1_exit219_S0: begin
        /* exec_result135 <= c2004 ? 0 : c2005 ? 0 : c2006 ? 1 : 'bz; */
        /* lit0_ip4 <= c2004 ? lit0_ip3 : c2005 ? lit0_ip2 : c2006 ? lit0_ip2 : 'bz; */
        /* lit0_phase6 <= c2004 ? 1 : c2005 ? 2 : c2006 ? 0 : 'bz; */
        /* stack0_pos4 <= c2004 ? stack0_pos2 : c2005 ? stack0_pos2 : c2006 ? stack0_pos3 : 'bz; */
        /* stack0_second4 <= c2004 ? stack0_second2 : c2005 ? stack0_second2 : c2006 ? stack0_top2 : 'bz; */
        /* stack0_top4 <= c2004 ? stack0_top2 : c2005 ? stack0_top2 : c2006 ? mem_data : 'bz; */
        retro_main_state <= retro_main_L1_b178_S0;
      end
      retro_main_L1_ifelse311_S5: begin
        _stack_addr <= t842_inl2_inl33;
        _stack_we <= 0;
        _stack_req <= 1;
        /* stack0_pos9 <= (stack0_pos2 - 1); */
        /* t842_inl2_inl33 <= (stack0_pos9 - 2); */
        retro_main_state <= retro_main_L1_ifelse311_S6;
      end
      retro_main_L1_ifelse311_S6: begin
        /*wait for output of _stack*/
        retro_main_state <= retro_main_L1_ifelse311_S7;
      end
      retro_main_L1_ifelse311_S7: begin
        stack0_second10 <= _stack_q;
        _stack_req <= 0;
        retro_main_state <= retro_main_L1_exit310_S0;
      end
      retro_main_L1_exit322_S0: begin
        /* c3404 <= (((c3346 && c882_inl34) || (c3346 && c1038_inl34)) || (c3346 && c1039_inl34)); */
        /* exec_result346 <= c2016 ? 0 : c2017 ? 0 : c2018 ? 0 : c2019 ? 1 : 'bz; */
        /* jump0_ip5 <= c2016 ? jump0_ip3 : c2017 ? jump0_ip2 : c2018 ? jump0_ip4 : c2019 ? jump0_ip2 : 'bz; */
        /* jump0_phase7 <= c2016 ? 1 : c2017 ? 2 : c2018 ? 3 : c2019 ? 0 : 'bz; */
        retro_main_state <= retro_main_L1_b178_S0;
      end
      retro_main_L1_b564_S0: begin
        /* t2771 <= c2126 ? 0 : c2127 ? 1 : 'bz; */
        /* t2774 <= c2126 ? 2 : c2127 ? 0 : 'bz; */
        retro_main_state <= retro_main_L1_exit333_S0;
      end
      retro_main_L1_b565_S0: begin
        /* t2778 <= c2128 ? 0 : c2129 ? 1 : 'bz; */
        /* t2781 <= c2128 ? 2 : c2129 ? 0 : 'bz; */
        retro_main_state <= retro_main_L1_exit350_S0;
      end
      retro_main_L1_b566_S0: begin
        /* t2785 <= c2130 ? 0 : c2131 ? 1 : 'bz; */
        /* t2788 <= c2130 ? 2 : c2131 ? 0 : 'bz; */
        retro_main_state <= retro_main_L1_exit367_S0;
      end
      retro_main_L1_b567_S0: begin
        /* t2792 <= c2132 ? 0 : c2133 ? 1 : 'bz; */
        /* t2795 <= c2132 ? 2 : c2133 ? 0 : 'bz; */
        retro_main_state <= retro_main_L1_exit384_S0;
      end
      retro_main_L1_exit397_S0: begin
        /* exec_result396 <= c2037 ? 0 : c2038 ? 0 : c2039 ? 0 : c2040 ? 1 : 'bz; */
        /* point0_ip5 <= c2037 ? stack0_top2 : c2038 ? point0_ip2 : c2039 ? point0_ip_saved2 : c2040 ? point0_ip2 : 'bz; */
        /* point0_ip_saved4 <= c2037 ? ip2 : c2038 ? point0_ip_saved2 : c2039 ? point0_ip_saved2 : c2040 ? point0_ip_saved2 : 'bz; */
        /* point0_phase7 <= c2037 ? 1 : c2038 ? 2 : c2039 ? 3 : c2040 ? 0 : 'bz; */
        /* stack0_top26 <= c2037 ? stack0_top2 : c2038 ? stack0_top2 : c2039 ? mem_data : c2040 ? stack0_top2 : 'bz; */
        retro_main_state <= retro_main_L1_b178_S0;
      end
      retro_main_L1_exit412_S0: begin
        /* exec_result404 <= c2041 ? 0 : c2042 ? 1 : 'bz; */
        /* stack0_pos25 <= c2041 ? stack0_pos23 : c2042 ? stack0_pos24 : 'bz; */
        /* stack0_second26 <= c2041 ? stack0_second24 : c2042 ? stack0_second25 : 'bz; */
        /* write_point0_addr4 <= c2041 ? stack0_top2 : c2042 ? write_point0_addr2 : 'bz; */
        /* write_point0_data4 <= c2041 ? write_point0_data2 : c2042 ? stack0_top2 : 'bz; */
        /* write_point0_ip4 <= c2041 ? ip2 : c2042 ? write_point0_ip2 : 'bz; */
        /* write_point0_phase5 <= c2041 ? 1 : c2042 ? 0 : 'bz; */
        /* c924 <= (exec_result404 != 0); */
        /* c2146 <= ((c2041 || c2042) && c924); */
        retro_main_state <= retro_main_L1_b568_S0;
      end
      retro_main_L1_ifthen479_S6: begin
        _address_addr <= t842_inl2_inl54;
        _address_we <= 0;
        _address_req <= 1;
        _stack_addr <= t842_inl1_inl54;
        _stack_we <= 0;
        _stack_req <= 1;
        /* stack0_pos34 <= (stack0_pos2 - 1); */
        /* address0_pos6 <= (address0_pos2 - 1); */
        /* t842_inl1_inl54 <= (stack0_pos34 - 2); */
        /* t842_inl2_inl54 <= (address0_pos6 - 2); */
        retro_main_state <= retro_main_L1_ifthen479_S7;
      end
      retro_main_L1_ifthen479_S7: begin
        /*wait for output of _address*/
        /*wait for output of _stack*/
        retro_main_state <= retro_main_L1_ifthen479_S8;
      end
      retro_main_L1_ifthen479_S8: begin
        address0_second6 <= _address_q;
        _address_req <= 0;
        stack0_second36 <= _stack_q;
        _stack_req <= 0;
        retro_main_state <= retro_main_L1_exit488_S0;
      end
      retro_main_L1_ifthen493_S1: begin
        array1010[1] <= 0;
        retro_main_state <= retro_main_L1_ifthen493_S2;
      end
      retro_main_L1_ifthen493_S2: begin
        t932_inl55 <= array1010[1];
        retro_main_state <= retro_main_L1_ifthen493_S3;
      end
      retro_main_L1_ifthen493_S3: begin
        /* c933_inl55 <= (t932_inl55 == 13); */
        /* c2120 <= (c2093 && c933_inl55); */
        if (c933_inl55) begin
          array1010[1] <= 10;
          /* c3408 <= (c3407 && c933_inl55); */
          retro_main_state <= retro_main_L1_b497_S0;
        end else begin
          t934_inl55 <= array1010[2];
          /* c3409 <= (c3401 && !c930_inl55); */
          /* c2139 <= (c2060 && !c930_inl55); */
          /* c3410 <= (c3407 && !c933_inl55); */
          /* c2140 <= (c2093 && !c933_inl55); */
          retro_main_state <= retro_main_L1_b497_S1;
        end
      end
      retro_main_L1_exit310_S0: begin
        exec_result336 <= c2124 ? exec_result336 : c2125 ? 1 : c2013 ? 0 : c2014 ? 0 : c2015 ? 1 : 'bz;
        /* loop0_ip5 <= c2124 ? loop0_ip3 : c2125 ? loop0_ip3 : c2013 ? loop0_ip2 : c2014 ? loop0_ip4 : c2015 ? loop0_ip2 : 'bz; */
        /* loop0_phase8 <= c2124 ? 1 : c2125 ? 0 : c2013 ? 2 : c2014 ? 3 : c2015 ? 0 : 'bz; */
        /* stack0_pos10 <= c2124 ? stack0_pos2 : c2125 ? stack0_pos9 : c2013 ? stack0_pos2 : c2014 ? stack0_pos2 : c2015 ? stack0_pos2 : 'bz; */
        /* stack0_second11 <= c2124 ? stack0_second2 : c2125 ? stack0_second10 : c2013 ? stack0_second2 : c2014 ? stack0_second2 : c2015 ? stack0_second2 : 'bz; */
        /* stack0_top12 <= c2124 ? stack0_top10 : c2125 ? stack0_second2 : c2013 ? stack0_top2 : c2014 ? stack0_top2 : c2015 ? stack0_top2 : 'bz; */
        retro_main_state <= retro_main_L1_b178_S0;
      end
      retro_main_L1_exit333_S0: begin
        /* jump_ge0_a4 <= c2021 ? stack0_top2 : c2022 ? jump_ge0_a2 : c2023 ? jump_ge0_a2 : c2024 ? jump_ge0_a2 : 'bz; */
        /* jump_ge0_ip5 <= c2021 ? jump_ge0_ip3 : c2022 ? jump_ge0_ip2 : c2023 ? jump_ge0_ip4 : c2024 ? jump_ge0_ip2 : 'bz; */
        /* stack0_pos13 <= c2021 ? stack0_pos11 : c2022 ? stack0_pos12 : c2023 ? stack0_pos2 : c2024 ? stack0_pos2 : 'bz; */
        /* stack0_second14 <= c2021 ? stack0_second12 : c2022 ? stack0_second13 : c2023 ? stack0_second2 : c2024 ? stack0_second2 : 'bz; */
        /* stack0_top15 <= c2021 ? stack0_second2 : c2022 ? stack0_second2 : c2023 ? stack0_top2 : c2024 ? stack0_top2 : 'bz; */
        /* exec_result357 <= c2021 ? 0 : c2022 ? t2771 : c2023 ? 0 : c2024 ? 1 : 'bz; */
        /* jump_ge0_phase8 <= c2021 ? 1 : c2022 ? t2774 : c2023 ? 3 : c2024 ? 0 : 'bz; */
        retro_main_state <= retro_main_L1_b178_S0;
      end
      retro_main_L1_exit350_S0: begin
        /* jump_le0_a4 <= c2025 ? stack0_top2 : c2026 ? jump_le0_a2 : c2027 ? jump_le0_a2 : c2028 ? jump_le0_a2 : 'bz; */
        /* jump_le0_ip5 <= c2025 ? jump_le0_ip3 : c2026 ? jump_le0_ip2 : c2027 ? jump_le0_ip4 : c2028 ? jump_le0_ip2 : 'bz; */
        /* stack0_pos16 <= c2025 ? stack0_pos14 : c2026 ? stack0_pos15 : c2027 ? stack0_pos2 : c2028 ? stack0_pos2 : 'bz; */
        /* stack0_second17 <= c2025 ? stack0_second15 : c2026 ? stack0_second16 : c2027 ? stack0_second2 : c2028 ? stack0_second2 : 'bz; */
        /* stack0_top18 <= c2025 ? stack0_second2 : c2026 ? stack0_second2 : c2027 ? stack0_top2 : c2028 ? stack0_top2 : 'bz; */
        /* exec_result367 <= c2025 ? 0 : c2026 ? t2778 : c2027 ? 0 : c2028 ? 1 : 'bz; */
        /* jump_le0_phase8 <= c2025 ? 1 : c2026 ? t2781 : c2027 ? 3 : c2028 ? 0 : 'bz; */
        retro_main_state <= retro_main_L1_b178_S0;
      end
      retro_main_L1_exit367_S0: begin
        /* jump_ne0_a4 <= c2029 ? stack0_top2 : c2030 ? jump_ne0_a2 : c2031 ? jump_ne0_a2 : c2032 ? jump_ne0_a2 : 'bz; */
        /* jump_ne0_ip5 <= c2029 ? jump_ne0_ip3 : c2030 ? jump_ne0_ip2 : c2031 ? jump_ne0_ip4 : c2032 ? jump_ne0_ip2 : 'bz; */
        /* stack0_pos19 <= c2029 ? stack0_pos17 : c2030 ? stack0_pos18 : c2031 ? stack0_pos2 : c2032 ? stack0_pos2 : 'bz; */
        /* stack0_second20 <= c2029 ? stack0_second18 : c2030 ? stack0_second19 : c2031 ? stack0_second2 : c2032 ? stack0_second2 : 'bz; */
        /* stack0_top21 <= c2029 ? stack0_second2 : c2030 ? stack0_second2 : c2031 ? stack0_top2 : c2032 ? stack0_top2 : 'bz; */
        /* exec_result377 <= c2029 ? 0 : c2030 ? t2785 : c2031 ? 0 : c2032 ? 1 : 'bz; */
        /* jump_ne0_phase8 <= c2029 ? 1 : c2030 ? t2788 : c2031 ? 3 : c2032 ? 0 : 'bz; */
        retro_main_state <= retro_main_L1_b178_S0;
      end
      retro_main_L1_exit384_S0: begin
        /* jump_eq0_a4 <= c2033 ? stack0_top2 : c2034 ? jump_eq0_a2 : c2035 ? jump_eq0_a2 : c2036 ? jump_eq0_a2 : 'bz; */
        /* jump_eq0_ip5 <= c2033 ? jump_eq0_ip3 : c2034 ? jump_eq0_ip2 : c2035 ? jump_eq0_ip4 : c2036 ? jump_eq0_ip2 : 'bz; */
        /* stack0_pos22 <= c2033 ? stack0_pos20 : c2034 ? stack0_pos21 : c2035 ? stack0_pos2 : c2036 ? stack0_pos2 : 'bz; */
        /* stack0_second23 <= c2033 ? stack0_second21 : c2034 ? stack0_second22 : c2035 ? stack0_second2 : c2036 ? stack0_second2 : 'bz; */
        /* stack0_top24 <= c2033 ? stack0_second2 : c2034 ? stack0_second2 : c2035 ? stack0_top2 : c2036 ? stack0_top2 : 'bz; */
        /* exec_result387 <= c2033 ? 0 : c2034 ? t2792 : c2035 ? 0 : c2036 ? 1 : 'bz; */
        /* jump_eq0_phase8 <= c2033 ? 1 : c2034 ? t2795 : c2035 ? 3 : c2036 ? 0 : 'bz; */
        retro_main_state <= retro_main_L1_b178_S0;
      end
      retro_main_L1_b568_S0: begin
        /* t2829 <= c2146 ? 1 : ((c2041 || c2042) && !c924) ? wr_flag2 : 'bz; */
        /* t2830 <= c2146 ? write_point0_addr4 : ((c2041 || c2042) && !c924) ? wr_mem_addr2 : 'bz; */
        /* t2831 <= c2146 ? write_point0_data4 : ((c2041 || c2042) && !c924) ? wr_mem_data2 : 'bz; */
        retro_main_state <= retro_main_L1_b178_S0;
      end
      retro_main_L1_exit488_S0: begin
        /* address0_pos7 <= c2090 ? address0_pos6 : c2091 ? address0_pos2 : c2055 ? address0_pos2 : 'bz; */
        /* address0_second7 <= c2090 ? address0_second6 : c2091 ? address0_second2 : c2055 ? address0_second2 : 'bz; */
        /* address0_top7 <= c2090 ? address0_second2 : c2091 ? address0_top2 : c2055 ? address0_top2 : 'bz; */
        /* exec_result545 <= c2090 ? 0 : c2091 ? 1 : c2055 ? 1 : 'bz; */
        /* stack0_pos35 <= c2090 ? stack0_pos34 : c2091 ? stack0_pos2 : c2055 ? stack0_pos2 : 'bz; */
        /* stack0_second37 <= c2090 ? stack0_second36 : c2091 ? stack0_second2 : c2055 ? stack0_second2 : 'bz; */
        /* stack0_top48 <= c2090 ? stack0_second2 : c2091 ? stack0_top2 : c2055 ? stack0_top2 : 'bz; */
        /* zero_pop_return0_ip5 <= c2090 ? address0_top2 : c2091 ? ip2 : c2055 ? zero_pop_return0_ip2 : 'bz; */
        /* zero_pop_return0_phase5 <= c2090 ? 1 : c2091 ? zero_pop_return0_phase2 : c2055 ? 0 : 'bz; */
        retro_main_state <= retro_main_L1_b178_S0;
      end
      retro_main_L1_b497_S0: begin
        t934_inl55 <= array1010[2];
        /* c3409 <= (c3401 && !c930_inl55); */
        /* c2139 <= (c2060 && !c930_inl55); */
        /* c3410 <= (c3407 && !c933_inl55); */
        /* c2140 <= (c2093 && !c933_inl55); */
        retro_main_state <= retro_main_L1_b497_S1;
      end
      retro_main_L1_b497_S1: begin
        /* c935_inl55 <= (t934_inl55 == 1); */
        if (c935_inl55) begin
          /* c936_inl55 <= (stack0_top2 > 0); */
          /* c937_inl55 <= (stack0_top2 < 128); */
          /* c938_inl55 <= (c936_inl55 && c937_inl55); */
          /* c3411 <= (((c3409 || c3410) || c3408) && c935_inl55); */
          /* c2148 <= (((c2139 || c2140) || c2120) && c935_inl55); */
          if (c938_inl55) begin
            /* c939_inl55 <= (stack0_top2 == 8); */
            /* c3412 <= (c3411 && c938_inl55); */
            /* c2151 <= (c2148 && c938_inl55); */
            if (c939_inl55) begin
              /* c3414 <= (c3412 && c939_inl55); */
              /* c2155 <= (c2151 && c939_inl55); */
              retro_main_state <= retro_main_L1_ifthen500_S6;
            end else begin
              /* c3415 <= (c3412 && !c939_inl55); */
              /* c2156 <= (c2151 && !c939_inl55); */
              retro_main_state <= retro_main_L1_ifelse551_S6;
            end
          end else begin
            /* c3413 <= (c3411 && !c938_inl55); */
            /* c2152 <= (c2148 && !c938_inl55); */
            retro_main_state <= retro_main_L1_ifelse558_S6;
          end
        end else begin
          t941_inl55 <= array1010[4];
          /* c3416 <= (((c3409 || c3410) || c3408) && !c935_inl55); */
          /* c2166 <= (((c2139 || c2140) || c2120) && !c935_inl55); */
          /* c3417 <= ((c3413 || c3414) || c3415); */
          /* stack0_top58 <= ((c2152 || c2155) || c2156) ? stack0_second2 : (((c2139 || c2140) || c2120) && !c935_inl55) ? stack0_top2 : 'bz; */
          /* c2167 <= ((c2152 || c2155) || c2156); */
          /* stack0_pos42 <= ((c2152 || c2155) || c2156) ? stack0_pos41 : (((c2139 || c2140) || c2120) && !c935_inl55) ? stack0_pos2 : 'bz; */
          /* stack0_second44 <= ((c2152 || c2155) || c2156) ? stack0_second43 : (((c2139 || c2140) || c2120) && !c935_inl55) ? stack0_second2 : 'bz; */
          retro_main_state <= retro_main_L1_b514_S1;
        end
      end
      retro_main_L1_ifelse558_S6: begin
        _stack_addr <= t842_inl4_inl55;
        _stack_we <= 0;
        _stack_req <= 1;
        /* stack0_pos40 <= (stack0_pos2 - 1); */
        /* t842_inl4_inl55 <= (stack0_pos40 - 2); */
        retro_main_state <= retro_main_L1_ifelse558_S7;
      end
      retro_main_L1_ifelse558_S7: begin
        /*wait for output of _stack*/
        retro_main_state <= retro_main_L1_ifelse558_S8;
      end
      retro_main_L1_ifelse558_S8: begin
        stack0_second42 <= _stack_q;
        _stack_req <= 0;
        retro_main_state <= retro_main_L1_b511_S0;
      end
      retro_main_L1_ifthen500_S6: begin
        _stack_addr <= t842_inl2_inl55;
        _stack_we <= 0;
        _stack_req <= 1;
        /* stack0_pos38 <= (stack0_pos2 - 1); */
        /* t842_inl2_inl55 <= (stack0_pos38 - 2); */
        retro_main_state <= retro_main_L1_ifthen500_S7;
      end
      retro_main_L1_ifthen500_S7: begin
        /*wait for output of _stack*/
        retro_main_state <= retro_main_L1_ifthen500_S8;
      end
      retro_main_L1_ifthen500_S8: begin
        stack0_second40 <= _stack_q;
        _stack_req <= 0;
        retro_main_state <= retro_main_L1_ifthen500_S9;
      end
      retro_main_L1_ifthen500_S9: begin
        $display("%1d", stack0_top2);
        retro_main_state <= retro_main_L1_ifthen500_S10;
      end
      retro_main_L1_ifthen500_S10: begin
        $display("%1d", 32);
        retro_main_state <= retro_main_L1_ifthen500_S11;
      end
      retro_main_L1_ifthen500_S11: begin
        $display("%1d", 8);
        retro_main_state <= retro_main_L1_b511_S0;
      end
      retro_main_L1_ifelse551_S6: begin
        _stack_addr <= t842_inl3_inl55;
        _stack_we <= 0;
        _stack_req <= 1;
        /* stack0_pos39 <= (stack0_pos2 - 1); */
        /* t842_inl3_inl55 <= (stack0_pos39 - 2); */
        retro_main_state <= retro_main_L1_ifelse551_S7;
      end
      retro_main_L1_ifelse551_S7: begin
        /*wait for output of _stack*/
        retro_main_state <= retro_main_L1_ifelse551_S8;
      end
      retro_main_L1_ifelse551_S8: begin
        stack0_second41 <= _stack_q;
        _stack_req <= 0;
        retro_main_state <= retro_main_L1_ifelse551_S9;
      end
      retro_main_L1_ifelse551_S9: begin
        $display("%1d", stack0_top2);
        retro_main_state <= retro_main_L1_b511_S0;
      end
      retro_main_L1_b511_S0: begin
        array1010[2] <= 0;
        /* stack0_pos41 <= c2155 ? stack0_pos38 : c2156 ? stack0_pos39 : c2152 ? stack0_pos40 : 'bz; */
        /* stack0_second43 <= c2155 ? stack0_second40 : c2156 ? stack0_second41 : c2152 ? stack0_second42 : 'bz; */
        retro_main_state <= retro_main_L1_b514_S0;
      end
      retro_main_L1_b514_S0: begin
        t941_inl55 <= array1010[4];
        /* c3416 <= (((c3409 || c3410) || c3408) && !c935_inl55); */
        /* c2166 <= (((c2139 || c2140) || c2120) && !c935_inl55); */
        /* c3417 <= ((c3413 || c3414) || c3415); */
        /* stack0_top58 <= ((c2152 || c2155) || c2156) ? stack0_second2 : (((c2139 || c2140) || c2120) && !c935_inl55) ? stack0_top2 : 'bz; */
        /* c2167 <= ((c2152 || c2155) || c2156); */
        /* stack0_pos42 <= ((c2152 || c2155) || c2156) ? stack0_pos41 : (((c2139 || c2140) || c2120) && !c935_inl55) ? stack0_pos2 : 'bz; */
        /* stack0_second44 <= ((c2152 || c2155) || c2156) ? stack0_second43 : (((c2139 || c2140) || c2120) && !c935_inl55) ? stack0_second2 : 'bz; */
        retro_main_state <= retro_main_L1_b514_S1;
      end
      retro_main_L1_b514_S1: begin
        /* c942_inl55 <= (t941_inl55 == 1); */
        /* c2168 <= ((c2166 || c2167) && c942_inl55); */
        if (c942_inl55) begin
          array1010[4] <= 0;
          /* c3418 <= ((c3416 || c3417) && c942_inl55); */
          retro_main_state <= retro_main_L1_b516_S0;
        end else begin
          t943_inl55 <= array1010[4];
          /* c3419 <= ((c3416 || c3417) && !c942_inl55); */
          /* c2169 <= ((c2166 || c2167) && !c942_inl55); */
          retro_main_state <= retro_main_L1_b516_S1;
        end
      end
      retro_main_L1_b516_S0: begin
        t943_inl55 <= array1010[4];
        /* c3419 <= ((c3416 || c3417) && !c942_inl55); */
        /* c2169 <= ((c2166 || c2167) && !c942_inl55); */
        retro_main_state <= retro_main_L1_b516_S1;
      end
      retro_main_L1_b516_S1: begin
        /* c944_inl55 <= (t943_inl55 == 2); */
        /* c2170 <= ((c2169 || c2168) && c944_inl55); */
        if (c944_inl55) begin
          array1010[4] <= 0;
          /* c3420 <= ((c3419 || c3418) && c944_inl55); */
          retro_main_state <= retro_main_L1_b518_S0;
        end else begin
          t945_inl55 <= array1010[4];
          t947_inl55 <= array1010[4];
          t949_inl55 <= array1010[4];
          t951_inl55 <= array1010[4];
          t953_inl55 <= array1010[4];
          t955_inl55 <= array1010[4];
          t957_inl55 <= array1010[4];
          /* c3421 <= ((c3419 || c3418) && !c944_inl55); */
          /* c2171 <= ((c2169 || c2168) && !c944_inl55); */
          retro_main_state <= retro_main_L1_b518_S1;
        end
      end
      retro_main_L1_b518_S0: begin
        t945_inl55 <= array1010[4];
        t947_inl55 <= array1010[4];
        t949_inl55 <= array1010[4];
        t951_inl55 <= array1010[4];
        t953_inl55 <= array1010[4];
        t955_inl55 <= array1010[4];
        t957_inl55 <= array1010[4];
        /* c3421 <= ((c3419 || c3418) && !c944_inl55); */
        /* c2171 <= ((c2169 || c2168) && !c944_inl55); */
        retro_main_state <= retro_main_L1_b518_S1;
      end
      retro_main_L1_b518_S1: begin
        /* c946_inl55 <= (t945_inl55 == -1); */
        /* c948_inl55 <= (t947_inl55 == -2); */
        /* c950_inl55 <= (t949_inl55 == -3); */
        /* c952_inl55 <= (t951_inl55 == -4); */
        /* c954_inl55 <= (t953_inl55 == -5); */
        /* c956_inl55 <= (t955_inl55 == -6); */
        /* c958_inl55 <= (t957_inl55 == -7); */
        /* c1072_inl55 <= (!c946_inl55 && c948_inl55); */
        /* c1073_inl55 <= ((!c946_inl55 && !c948_inl55) && c950_inl55); */
        /* c1074_inl55 <= (((!c946_inl55 && !c948_inl55) && !c950_inl55) && c952_inl55); */
        /* c1075_inl55 <= ((((!c946_inl55 && !c948_inl55) && !c950_inl55) && !c952_inl55) && c954_inl55); */
        /* c1076_inl55 <= (((((!c946_inl55 && !c948_inl55) && !c950_inl55) && !c952_inl55) && !c954_inl55) && c956_inl55); */
        /* c1077_inl55 <= ((((((!c946_inl55 && !c948_inl55) && !c950_inl55) && !c952_inl55) && !c954_inl55) && !c956_inl55) && c958_inl55); */
        /* c1078_inl55 <= ((((((!c946_inl55 && !c948_inl55) && !c950_inl55) && !c952_inl55) && !c954_inl55) && !c956_inl55) && !c958_inl55); */
        /* c2172 <= ((c2171 || c2170) && c946_inl55); */
        /* c2173 <= ((c2171 || c2170) && c1072_inl55); */
        /* c2174 <= ((c2171 || c2170) && c1073_inl55); */
        /* c2175 <= ((c2171 || c2170) && c1074_inl55); */
        /* c2176 <= ((c2171 || c2170) && c1075_inl55); */
        /* c2177 <= ((c2171 || c2170) && c1076_inl55); */
        /* c2178 <= ((c2171 || c2170) && c1077_inl55); */
        if (c946_inl55) begin
          array1010[4] <= 0;
          /* c3422 <= ((c3421 || c3420) && c946_inl55); */
          retro_main_state <= retro_main_L1_b520_S0;
        end else if (c1072_inl55) begin
          array1010[4] <= 0;
          /* c3423 <= ((c3421 || c3420) && c1072_inl55); */
          retro_main_state <= retro_main_L1_b520_S0;
        end else if (c1073_inl55) begin
          array1010[4] <= 1;
          /* c3424 <= ((c3421 || c3420) && c1073_inl55); */
          retro_main_state <= retro_main_L1_b520_S0;
        end else if (c1074_inl55) begin
          array1010[4] <= 0;
          /* c3425 <= ((c3421 || c3420) && c1074_inl55); */
          retro_main_state <= retro_main_L1_b520_S0;
        end else if (c1075_inl55) begin
          array1010[4] <= 0;
          /* c3426 <= ((c3421 || c3420) && c1075_inl55); */
          retro_main_state <= retro_main_L1_b520_S0;
        end else if (c1076_inl55) begin
          array1010[4] <= 0;
          /* c3427 <= ((c3421 || c3420) && c1076_inl55); */
          retro_main_state <= retro_main_L1_b520_S0;
        end else if (c1077_inl55) begin
          array1010[4] <= 0;
          /* c3428 <= ((c3421 || c3420) && c1077_inl55); */
          retro_main_state <= retro_main_L1_b520_S0;
        end else if (c1078_inl55) begin
          t959_inl55 <= array1010[4];
          /* c3429 <= ((c3421 || c3420) && c1078_inl55); */
          /* c2179 <= ((c2171 || c2170) && c1078_inl55); */
          retro_main_state <= retro_main_L1_b520_S1;
        end
      end
      retro_main_L1_b520_S0: begin
        t959_inl55 <= array1010[4];
        /* c3429 <= ((c3421 || c3420) && c1078_inl55); */
        /* c2179 <= ((c2171 || c2170) && c1078_inl55); */
        retro_main_state <= retro_main_L1_b520_S1;
      end
      retro_main_L1_b520_S1: begin
        /* c960_inl55 <= (t959_inl55 == -8); */
        /* c2180 <= ((((((((c2179 || c2177) || c2176) || c2175) || c2174) || c2173) || c2172) || c2178) && c960_inl55); */
        if (c960_inl55) begin
          array1010[4] <= 0;
          /* c3430 <= ((((((((c3429 || c3427) || c3426) || c3425) || c3424) || c3423) || c3422) || c3428) && c960_inl55); */
          retro_main_state <= retro_main_L1_b522_S0;
        end else begin
          t961_inl55 <= array1010[5];
          t963_inl55 <= array1010[5];
          t965_inl55 <= array1010[5];
          t967_inl55 <= array1010[5];
          t969_inl55 <= array1010[5];
          t971_inl55 <= array1010[5];
          t973_inl55 <= array1010[5];
          t975_inl55 <= array1010[5];
          t977_inl55 <= array1010[5];
          t979_inl55 <= array1010[5];
          t981_inl55 <= array1010[5];
          t983_inl55 <= array1010[5];
          t985_inl55 <= array1010[5];
          t987_inl55 <= array1010[5];
          t989_inl55 <= array1010[5];
          /* c3431 <= ((((((((c3429 || c3427) || c3426) || c3425) || c3424) || c3423) || c3422) || c3428) && !c960_inl55); */
          /* c2181 <= ((((((((c2179 || c2177) || c2176) || c2175) || c2174) || c2173) || c2172) || c2178) && !c960_inl55); */
          retro_main_state <= retro_main_L1_b522_S1;
        end
      end
      retro_main_L1_b522_S0: begin
        t961_inl55 <= array1010[5];
        t963_inl55 <= array1010[5];
        t965_inl55 <= array1010[5];
        t967_inl55 <= array1010[5];
        t969_inl55 <= array1010[5];
        t971_inl55 <= array1010[5];
        t973_inl55 <= array1010[5];
        t975_inl55 <= array1010[5];
        t977_inl55 <= array1010[5];
        t979_inl55 <= array1010[5];
        t981_inl55 <= array1010[5];
        t983_inl55 <= array1010[5];
        t985_inl55 <= array1010[5];
        t987_inl55 <= array1010[5];
        t989_inl55 <= array1010[5];
        /* c3431 <= ((((((((c3429 || c3427) || c3426) || c3425) || c3424) || c3423) || c3422) || c3428) && !c960_inl55); */
        /* c2181 <= ((((((((c2179 || c2177) || c2176) || c2175) || c2174) || c2173) || c2172) || c2178) && !c960_inl55); */
        retro_main_state <= retro_main_L1_b522_S1;
      end
      retro_main_L1_b522_S1: begin
        /* c962_inl55 <= (t961_inl55 == -1); */
        /* c964_inl55 <= (t963_inl55 == -2); */
        /* c966_inl55 <= (t965_inl55 == -3); */
        /* c968_inl55 <= (t967_inl55 == -4); */
        /* c970_inl55 <= (t969_inl55 == -5); */
        /* c972_inl55 <= (t971_inl55 == -6); */
        /* c974_inl55 <= (t973_inl55 == -7); */
        /* c976_inl55 <= (t975_inl55 == -8); */
        /* c978_inl55 <= (t977_inl55 == -9); */
        /* c980_inl55 <= (t979_inl55 == -10); */
        /* c982_inl55 <= (t981_inl55 == -11); */
        /* c984_inl55 <= (t983_inl55 == -12); */
        /* c986_inl55 <= (t985_inl55 == -13); */
        /* c988_inl55 <= (t987_inl55 == -14); */
        /* c990_inl55 <= (t989_inl55 == -15); */
        /* c1079_inl55 <= (!c962_inl55 && c964_inl55); */
        /* c1080_inl55 <= ((!c962_inl55 && !c964_inl55) && c966_inl55); */
        /* c1081_inl55 <= (((!c962_inl55 && !c964_inl55) && !c966_inl55) && c968_inl55); */
        /* c1082_inl55 <= ((((!c962_inl55 && !c964_inl55) && !c966_inl55) && !c968_inl55) && c970_inl55); */
        /* c1083_inl55 <= (((((!c962_inl55 && !c964_inl55) && !c966_inl55) && !c968_inl55) && !c970_inl55) && c972_inl55); */
        /* c1084_inl55 <= ((((((!c962_inl55 && !c964_inl55) && !c966_inl55) && !c968_inl55) && !c970_inl55) && !c972_inl55) && c974_inl55); */
        /* c1085_inl55 <= (((((((!c962_inl55 && !c964_inl55) && !c966_inl55) && !c968_inl55) && !c970_inl55) && !c972_inl55) && !c974_inl55) && c976_inl55); */
        /* c1086_inl55 <= ((((((((!c962_inl55 && !c964_inl55) && !c966_inl55) && !c968_inl55) && !c970_inl55) && !c972_inl55) && !c974_inl55) && !c976_inl55) && c978_inl55); */
        /* c1087_inl55 <= (((((((((!c962_inl55 && !c964_inl55) && !c966_inl55) && !c968_inl55) && !c970_inl55) && !c972_inl55) && !c974_inl55) && !c976_inl55) && !c978_inl55) && c980_inl55); */
        /* c1088_inl55 <= ((((((((((!c962_inl55 && !c964_inl55) && !c966_inl55) && !c968_inl55) && !c970_inl55) && !c972_inl55) && !c974_inl55) && !c976_inl55) && !c978_inl55) && !c980_inl55) && c982_inl55); */
        /* c1089_inl55 <= (((((((((((!c962_inl55 && !c964_inl55) && !c966_inl55) && !c968_inl55) && !c970_inl55) && !c972_inl55) && !c974_inl55) && !c976_inl55) && !c978_inl55) && !c980_inl55) && !c982_inl55) && c984_inl55); */
        /* c1090_inl55 <= ((((((((((((!c962_inl55 && !c964_inl55) && !c966_inl55) && !c968_inl55) && !c970_inl55) && !c972_inl55) && !c974_inl55) && !c976_inl55) && !c978_inl55) && !c980_inl55) && !c982_inl55) && !c984_inl55) && c986_inl55); */
        /* c1091_inl55 <= (((((((((((((!c962_inl55 && !c964_inl55) && !c966_inl55) && !c968_inl55) && !c970_inl55) && !c972_inl55) && !c974_inl55) && !c976_inl55) && !c978_inl55) && !c980_inl55) && !c982_inl55) && !c984_inl55) && !c986_inl55) && c988_inl55); */
        /* c1092_inl55 <= ((((((((((((((!c962_inl55 && !c964_inl55) && !c966_inl55) && !c968_inl55) && !c970_inl55) && !c972_inl55) && !c974_inl55) && !c976_inl55) && !c978_inl55) && !c980_inl55) && !c982_inl55) && !c984_inl55) && !c986_inl55) && !c988_inl55) && c990_inl55); */
        /* c1093_inl55 <= ((((((((((((((!c962_inl55 && !c964_inl55) && !c966_inl55) && !c968_inl55) && !c970_inl55) && !c972_inl55) && !c974_inl55) && !c976_inl55) && !c978_inl55) && !c980_inl55) && !c982_inl55) && !c984_inl55) && !c986_inl55) && !c988_inl55) && !c990_inl55); */
        /* c2182 <= ((c2181 || c2180) && c962_inl55); */
        /* c2183 <= ((c2181 || c2180) && c1079_inl55); */
        /* c2184 <= ((c2181 || c2180) && c1080_inl55); */
        /* c2185 <= ((c2181 || c2180) && c1081_inl55); */
        /* c2186 <= ((c2181 || c2180) && c1082_inl55); */
        /* c2187 <= ((c2181 || c2180) && c1083_inl55); */
        /* c2188 <= ((c2181 || c2180) && c1084_inl55); */
        /* c2189 <= ((c2181 || c2180) && c1085_inl55); */
        /* c2190 <= ((c2181 || c2180) && c1086_inl55); */
        /* c2191 <= ((c2181 || c2180) && c1087_inl55); */
        /* c2192 <= ((c2181 || c2180) && c1088_inl55); */
        /* c2193 <= ((c2181 || c2180) && c1089_inl55); */
        /* c2194 <= ((c2181 || c2180) && c1090_inl55); */
        /* c2195 <= ((c2181 || c2180) && c1091_inl55); */
        /* c2196 <= ((c2181 || c2180) && c1092_inl55); */
        if (c962_inl55) begin
          array1010[5] <= 99999;
          /* c3432 <= ((c3431 || c3430) && c962_inl55); */
          retro_main_state <= retro_main_L1_b524_S0;
        end else if (c1079_inl55) begin
          array1010[5] <= 0;
          /* c3433 <= ((c3431 || c3430) && c1079_inl55); */
          retro_main_state <= retro_main_L1_b524_S0;
        end else if (c1080_inl55) begin
          array1010[5] <= 0;
          /* c3434 <= ((c3431 || c3430) && c1080_inl55); */
          retro_main_state <= retro_main_L1_b524_S0;
        end else if (c1081_inl55) begin
          array1010[5] <= 0;
          /* c3435 <= ((c3431 || c3430) && c1081_inl55); */
          retro_main_state <= retro_main_L1_b524_S0;
        end else if (c1082_inl55) begin
          array1010[5] <= 128;
          /* c3436 <= ((c3431 || c3430) && c1082_inl55); */
          retro_main_state <= retro_main_L1_b524_S0;
        end else if (c1083_inl55) begin
          array1010[5] <= 1024;
          /* c3437 <= ((c3431 || c3430) && c1083_inl55); */
          retro_main_state <= retro_main_L1_b524_S0;
        end else if (c1084_inl55) begin
          array1010[5] <= 0;
          /* c3438 <= ((c3431 || c3430) && c1084_inl55); */
          retro_main_state <= retro_main_L1_b524_S0;
        end else if (c1085_inl55) begin
          array1010[5] <= 0;
          /* c3439 <= ((c3431 || c3430) && c1085_inl55); */
          retro_main_state <= retro_main_L1_b524_S0;
        end else if (c1086_inl55) begin
          array1010[5] <= 0;
          /* c3440 <= ((c3431 || c3430) && c1086_inl55); */
          retro_main_state <= retro_main_L1_b524_S0;
        end else if (c1087_inl55) begin
          array1010[5] <= 0;
          /* c3441 <= ((c3431 || c3430) && c1087_inl55); */
          retro_main_state <= retro_main_L1_b524_S0;
        end else if (c1088_inl55) begin
          array1010[5] <= 0;
          /* c3442 <= ((c3431 || c3430) && c1088_inl55); */
          retro_main_state <= retro_main_L1_b524_S0;
        end else if (c1089_inl55) begin
          array1010[5] <= 0;
          /* c3443 <= ((c3431 || c3430) && c1089_inl55); */
          retro_main_state <= retro_main_L1_b524_S0;
        end else if (c1090_inl55) begin
          array1010[5] <= 32;
          /* c3444 <= ((c3431 || c3430) && c1090_inl55); */
          retro_main_state <= retro_main_L1_b524_S0;
        end else if (c1091_inl55) begin
          array1010[5] <= 0;
          /* c3445 <= ((c3431 || c3430) && c1091_inl55); */
          retro_main_state <= retro_main_L1_b524_S0;
        end else if (c1092_inl55) begin
          array1010[5] <= -1;
          /* c3446 <= ((c3431 || c3430) && c1092_inl55); */
          retro_main_state <= retro_main_L1_b524_S0;
        end else if (c1093_inl55) begin
          t991_inl55 <= array1010[8];
          /* c3447 <= ((c3431 || c3430) && c1093_inl55); */
          /* c2197 <= ((c2181 || c2180) && c1093_inl55); */
          /* ip_inl554 <= c2182 ? ip2 : c2183 ? ip2 : c2184 ? ip2 : c2185 ? ip2 : c2186 ? ip2 : c2187 ? ip2 : c2188 ? ip2 : c2189 ? ip2 : c2190 ? 268435455 : c2191 ? ip2 : c2192 ? ip2 : c2193 ? ip2 : c2194 ? ip2 : c2195 ? ip2 : c2196 ? ip2 : ((c2181 || c2180) && c1093_inl55) ? ip2 : 'bz; */
          retro_main_state <= retro_main_L1_b524_S1;
        end
      end
      retro_main_L1_b524_S0: begin
        t991_inl55 <= array1010[8];
        /* c3447 <= ((c3431 || c3430) && c1093_inl55); */
        /* c2197 <= ((c2181 || c2180) && c1093_inl55); */
        /* ip_inl554 <= c2182 ? ip2 : c2183 ? ip2 : c2184 ? ip2 : c2185 ? ip2 : c2186 ? ip2 : c2187 ? ip2 : c2188 ? ip2 : c2189 ? ip2 : c2190 ? 268435455 : c2191 ? ip2 : c2192 ? ip2 : c2193 ? ip2 : c2194 ? ip2 : c2195 ? ip2 : c2196 ? ip2 : ((c2181 || c2180) && c1093_inl55) ? ip2 : 'bz; */
        retro_main_state <= retro_main_L1_b524_S1;
      end
      retro_main_L1_b524_S1: begin
        /* c992_inl55 <= (t991_inl55 == 1); */
        /* c2198 <= ((((((((((((((((c2197 || c2185) || c2195) || c2189) || c2194) || c2193) || c2191) || c2192) || c2184) || c2187) || c2190) || c2183) || c2182) || c2196) || c2186) || c2188) && c992_inl55); */
        if (c992_inl55) begin
          array1010[8] <= 0;
          /* c3448 <= ((((((((((((((((c3447 || c3435) || c3445) || c3439) || c3444) || c3443) || c3441) || c3442) || c3434) || c3437) || c3440) || c3433) || c3432) || c3446) || c3436) || c3438) && c992_inl55); */
          retro_main_state <= retro_main_L1_b526_S0;
        end else begin
          /* c3449 <= ((((((((((((((((c3447 || c3435) || c3445) || c3439) || c3444) || c3443) || c3441) || c3442) || c3434) || c3437) || c3440) || c3433) || c3432) || c3446) || c3436) || c3438) && !c992_inl55); */
          /* c2199 <= ((((((((((((((((c2197 || c2185) || c2195) || c2189) || c2194) || c2193) || c2191) || c2192) || c2184) || c2187) || c2190) || c2183) || c2182) || c2196) || c2186) || c2188) && !c992_inl55); */
          retro_main_state <= retro_main_L1_b178_S0;
        end
      end
      retro_main_L1_b526_S0: begin
        /* c3449 <= ((((((((((((((((c3447 || c3435) || c3445) || c3439) || c3444) || c3443) || c3441) || c3442) || c3434) || c3437) || c3440) || c3433) || c3432) || c3446) || c3436) || c3438) && !c992_inl55); */
        /* c2199 <= ((((((((((((((((c2197 || c2185) || c2195) || c2189) || c2194) || c2193) || c2191) || c2192) || c2184) || c2187) || c2190) || c2183) || c2182) || c2196) || c2186) || c2188) && !c992_inl55); */
        retro_main_state <= retro_main_L1_b178_S0;
      end
      retro_main_L1_b178_S0: begin
        /* address0_pos9 <= (c1971 && c889) ? address0_pos2 : ((c2004 || c2005) || c2006) ? address0_pos2 : c1974 ? address0_pos2 : c1975 ? address0_pos2 : c1976 ? address0_pos2 : c1977 ? address0_pos3 : c1978 ? address0_pos4 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? address0_pos2 : (((c2019 || c2017) || c2018) || c2016) ? address0_pos2 : c1981 ? address0_pos5 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? address0_pos2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? address0_pos2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? address0_pos2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? address0_pos2 : (((c2038 || c2040) || c2037) || c2039) ? address0_pos2 : (c2041 || c2042) ? address0_pos2 : c1988 ? address0_pos2 : c1989 ? address0_pos2 : c1990 ? address0_pos2 : c1991 ? address0_pos2 : c1992 ? address0_pos2 : c1993 ? address0_pos2 : c1994 ? address0_pos2 : c1995 ? address0_pos2 : c1996 ? address0_pos2 : ((c2055 || c2091) || c2090) ? address0_pos7 : c1998 ? address0_pos2 : c1999 ? address0_pos2 : c2000 ? address0_pos2 : c2001 ? address0_pos2 : (c2199 || c2198) ? address0_pos2 : (c2002 && !c927) ? address0_pos2 : c1972 ? address0_pos8 : 'bz; */
        /* address0_second9 <= (c1971 && c889) ? address0_second2 : ((c2004 || c2005) || c2006) ? address0_second2 : c1974 ? address0_second2 : c1975 ? address0_second2 : c1976 ? address0_second2 : c1977 ? address0_top2 : c1978 ? address0_second4 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? address0_second2 : (((c2019 || c2017) || c2018) || c2016) ? address0_second2 : c1981 ? address0_second5 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? address0_second2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? address0_second2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? address0_second2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? address0_second2 : (((c2038 || c2040) || c2037) || c2039) ? address0_second2 : (c2041 || c2042) ? address0_second2 : c1988 ? address0_second2 : c1989 ? address0_second2 : c1990 ? address0_second2 : c1991 ? address0_second2 : c1992 ? address0_second2 : c1993 ? address0_second2 : c1994 ? address0_second2 : c1995 ? address0_second2 : c1996 ? address0_second2 : ((c2055 || c2091) || c2090) ? address0_second7 : c1998 ? address0_second2 : c1999 ? address0_second2 : c2000 ? address0_second2 : c2001 ? address0_second2 : (c2199 || c2198) ? address0_second2 : (c2002 && !c927) ? address0_second2 : c1972 ? address0_top2 : 'bz; */
        /* address0_top9 <= (c1971 && c889) ? address0_top2 : ((c2004 || c2005) || c2006) ? address0_top2 : c1974 ? address0_top2 : c1975 ? address0_top2 : c1976 ? address0_top2 : c1977 ? stack0_top2 : c1978 ? address0_second2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? address0_top2 : (((c2019 || c2017) || c2018) || c2016) ? address0_top2 : c1981 ? address0_second2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? address0_top2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? address0_top2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? address0_top2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? address0_top2 : (((c2038 || c2040) || c2037) || c2039) ? address0_top2 : (c2041 || c2042) ? address0_top2 : c1988 ? address0_top2 : c1989 ? address0_top2 : c1990 ? address0_top2 : c1991 ? address0_top2 : c1992 ? address0_top2 : c1993 ? address0_top2 : c1994 ? address0_top2 : c1995 ? address0_top2 : c1996 ? address0_top2 : ((c2055 || c2091) || c2090) ? address0_top7 : c1998 ? address0_top2 : c1999 ? address0_top2 : c2000 ? address0_top2 : c2001 ? address0_top2 : (c2199 || c2198) ? address0_top2 : (c2002 && !c927) ? address0_top2 : c1972 ? ip2 : 'bz; */
        /* done_flag13 <= (c1971 && c889) ? done_flag2 : ((c2004 || c2005) || c2006) ? exec_result135 : c1974 ? done_flag2 : c1975 ? done_flag2 : c1976 ? done_flag2 : c1977 ? done_flag2 : c1978 ? done_flag2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? exec_result336 : (((c2019 || c2017) || c2018) || c2016) ? exec_result346 : c1981 ? done_flag2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? exec_result357 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? exec_result367 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? exec_result377 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? exec_result387 : (((c2038 || c2040) || c2037) || c2039) ? exec_result396 : (c2041 || c2042) ? exec_result404 : c1988 ? done_flag2 : c1989 ? done_flag2 : c1990 ? done_flag2 : c1991 ? done_flag2 : c1992 ? done_flag2 : c1993 ? done_flag2 : c1994 ? done_flag2 : c1995 ? done_flag2 : c1996 ? done_flag2 : ((c2055 || c2091) || c2090) ? exec_result545 : c1998 ? done_flag2 : c1999 ? done_flag2 : c2000 ? done_flag2 : c2001 ? done_flag2 : (c2199 || c2198) ? done_flag2 : (c2002 && !c927) ? done_flag2 : c1972 ? done_flag2 : 'bz; */
        /* ip16 <= (c1971 && c889) ? ip2 : ((c2004 || c2005) || c2006) ? lit0_ip4 : c1974 ? ip2 : c1975 ? ip2 : c1976 ? ip2 : c1977 ? ip2 : c1978 ? ip2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? loop0_ip5 : (((c2019 || c2017) || c2018) || c2016) ? jump0_ip5 : c1981 ? address0_top2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? jump_ge0_ip5 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? jump_le0_ip5 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? jump_ne0_ip5 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? jump_eq0_ip5 : (((c2038 || c2040) || c2037) || c2039) ? point0_ip5 : (c2041 || c2042) ? write_point0_ip4 : c1988 ? ip2 : c1989 ? ip2 : c1990 ? ip2 : c1991 ? ip2 : c1992 ? ip2 : c1993 ? ip2 : c1994 ? ip2 : c1995 ? ip2 : c1996 ? ip2 : ((c2055 || c2091) || c2090) ? zero_pop_return0_ip5 : c1998 ? ip2 : c1999 ? ip2 : c2000 ? ip2 : c2001 ? ip2 : (c2199 || c2198) ? ip_inl554 : (c2002 && !c927) ? ip2 : c1972 ? ip15 : 'bz; */
        /* jump0_ip6 <= (c1971 && c889) ? jump0_ip2 : ((c2004 || c2005) || c2006) ? jump0_ip2 : c1974 ? jump0_ip2 : c1975 ? jump0_ip2 : c1976 ? jump0_ip2 : c1977 ? jump0_ip2 : c1978 ? jump0_ip2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? jump0_ip2 : (((c2019 || c2017) || c2018) || c2016) ? jump0_ip5 : c1981 ? jump0_ip2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? jump0_ip2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? jump0_ip2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? jump0_ip2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? jump0_ip2 : (((c2038 || c2040) || c2037) || c2039) ? jump0_ip2 : (c2041 || c2042) ? jump0_ip2 : c1988 ? jump0_ip2 : c1989 ? jump0_ip2 : c1990 ? jump0_ip2 : c1991 ? jump0_ip2 : c1992 ? jump0_ip2 : c1993 ? jump0_ip2 : c1994 ? jump0_ip2 : c1995 ? jump0_ip2 : c1996 ? jump0_ip2 : ((c2055 || c2091) || c2090) ? jump0_ip2 : c1998 ? jump0_ip2 : c1999 ? jump0_ip2 : c2000 ? jump0_ip2 : c2001 ? jump0_ip2 : (c2199 || c2198) ? jump0_ip2 : (c2002 && !c927) ? jump0_ip2 : c1972 ? jump0_ip2 : 'bz; */
        /* jump0_phase8 <= (c1971 && c889) ? jump0_phase2 : ((c2004 || c2005) || c2006) ? jump0_phase2 : c1974 ? jump0_phase2 : c1975 ? jump0_phase2 : c1976 ? jump0_phase2 : c1977 ? jump0_phase2 : c1978 ? jump0_phase2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? jump0_phase2 : (((c2019 || c2017) || c2018) || c2016) ? jump0_phase7 : c1981 ? jump0_phase2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? jump0_phase2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? jump0_phase2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? jump0_phase2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? jump0_phase2 : (((c2038 || c2040) || c2037) || c2039) ? jump0_phase2 : (c2041 || c2042) ? jump0_phase2 : c1988 ? jump0_phase2 : c1989 ? jump0_phase2 : c1990 ? jump0_phase2 : c1991 ? jump0_phase2 : c1992 ? jump0_phase2 : c1993 ? jump0_phase2 : c1994 ? jump0_phase2 : c1995 ? jump0_phase2 : c1996 ? jump0_phase2 : ((c2055 || c2091) || c2090) ? jump0_phase2 : c1998 ? jump0_phase2 : c1999 ? jump0_phase2 : c2000 ? jump0_phase2 : c2001 ? jump0_phase2 : (c2199 || c2198) ? jump0_phase2 : (c2002 && !c927) ? jump0_phase2 : c1972 ? jump0_phase2 : 'bz; */
        /* jump_eq0_a5 <= (c1971 && c889) ? jump_eq0_a2 : ((c2004 || c2005) || c2006) ? jump_eq0_a2 : c1974 ? jump_eq0_a2 : c1975 ? jump_eq0_a2 : c1976 ? jump_eq0_a2 : c1977 ? jump_eq0_a2 : c1978 ? jump_eq0_a2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? jump_eq0_a2 : (((c2019 || c2017) || c2018) || c2016) ? jump_eq0_a2 : c1981 ? jump_eq0_a2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? jump_eq0_a2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? jump_eq0_a2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? jump_eq0_a2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? jump_eq0_a4 : (((c2038 || c2040) || c2037) || c2039) ? jump_eq0_a2 : (c2041 || c2042) ? jump_eq0_a2 : c1988 ? jump_eq0_a2 : c1989 ? jump_eq0_a2 : c1990 ? jump_eq0_a2 : c1991 ? jump_eq0_a2 : c1992 ? jump_eq0_a2 : c1993 ? jump_eq0_a2 : c1994 ? jump_eq0_a2 : c1995 ? jump_eq0_a2 : c1996 ? jump_eq0_a2 : ((c2055 || c2091) || c2090) ? jump_eq0_a2 : c1998 ? jump_eq0_a2 : c1999 ? jump_eq0_a2 : c2000 ? jump_eq0_a2 : c2001 ? jump_eq0_a2 : (c2199 || c2198) ? jump_eq0_a2 : (c2002 && !c927) ? jump_eq0_a2 : c1972 ? jump_eq0_a2 : 'bz; */
        /* jump_eq0_ip6 <= (c1971 && c889) ? jump_eq0_ip2 : ((c2004 || c2005) || c2006) ? jump_eq0_ip2 : c1974 ? jump_eq0_ip2 : c1975 ? jump_eq0_ip2 : c1976 ? jump_eq0_ip2 : c1977 ? jump_eq0_ip2 : c1978 ? jump_eq0_ip2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? jump_eq0_ip2 : (((c2019 || c2017) || c2018) || c2016) ? jump_eq0_ip2 : c1981 ? jump_eq0_ip2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? jump_eq0_ip2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? jump_eq0_ip2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? jump_eq0_ip2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? jump_eq0_ip5 : (((c2038 || c2040) || c2037) || c2039) ? jump_eq0_ip2 : (c2041 || c2042) ? jump_eq0_ip2 : c1988 ? jump_eq0_ip2 : c1989 ? jump_eq0_ip2 : c1990 ? jump_eq0_ip2 : c1991 ? jump_eq0_ip2 : c1992 ? jump_eq0_ip2 : c1993 ? jump_eq0_ip2 : c1994 ? jump_eq0_ip2 : c1995 ? jump_eq0_ip2 : c1996 ? jump_eq0_ip2 : ((c2055 || c2091) || c2090) ? jump_eq0_ip2 : c1998 ? jump_eq0_ip2 : c1999 ? jump_eq0_ip2 : c2000 ? jump_eq0_ip2 : c2001 ? jump_eq0_ip2 : (c2199 || c2198) ? jump_eq0_ip2 : (c2002 && !c927) ? jump_eq0_ip2 : c1972 ? jump_eq0_ip2 : 'bz; */
        /* jump_eq0_phase9 <= (c1971 && c889) ? jump_eq0_phase2 : ((c2004 || c2005) || c2006) ? jump_eq0_phase2 : c1974 ? jump_eq0_phase2 : c1975 ? jump_eq0_phase2 : c1976 ? jump_eq0_phase2 : c1977 ? jump_eq0_phase2 : c1978 ? jump_eq0_phase2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? jump_eq0_phase2 : (((c2019 || c2017) || c2018) || c2016) ? jump_eq0_phase2 : c1981 ? jump_eq0_phase2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? jump_eq0_phase2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? jump_eq0_phase2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? jump_eq0_phase2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? jump_eq0_phase8 : (((c2038 || c2040) || c2037) || c2039) ? jump_eq0_phase2 : (c2041 || c2042) ? jump_eq0_phase2 : c1988 ? jump_eq0_phase2 : c1989 ? jump_eq0_phase2 : c1990 ? jump_eq0_phase2 : c1991 ? jump_eq0_phase2 : c1992 ? jump_eq0_phase2 : c1993 ? jump_eq0_phase2 : c1994 ? jump_eq0_phase2 : c1995 ? jump_eq0_phase2 : c1996 ? jump_eq0_phase2 : ((c2055 || c2091) || c2090) ? jump_eq0_phase2 : c1998 ? jump_eq0_phase2 : c1999 ? jump_eq0_phase2 : c2000 ? jump_eq0_phase2 : c2001 ? jump_eq0_phase2 : (c2199 || c2198) ? jump_eq0_phase2 : (c2002 && !c927) ? jump_eq0_phase2 : c1972 ? jump_eq0_phase2 : 'bz; */
        /* jump_ge0_a5 <= (c1971 && c889) ? jump_ge0_a2 : ((c2004 || c2005) || c2006) ? jump_ge0_a2 : c1974 ? jump_ge0_a2 : c1975 ? jump_ge0_a2 : c1976 ? jump_ge0_a2 : c1977 ? jump_ge0_a2 : c1978 ? jump_ge0_a2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? jump_ge0_a2 : (((c2019 || c2017) || c2018) || c2016) ? jump_ge0_a2 : c1981 ? jump_ge0_a2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? jump_ge0_a4 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? jump_ge0_a2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? jump_ge0_a2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? jump_ge0_a2 : (((c2038 || c2040) || c2037) || c2039) ? jump_ge0_a2 : (c2041 || c2042) ? jump_ge0_a2 : c1988 ? jump_ge0_a2 : c1989 ? jump_ge0_a2 : c1990 ? jump_ge0_a2 : c1991 ? jump_ge0_a2 : c1992 ? jump_ge0_a2 : c1993 ? jump_ge0_a2 : c1994 ? jump_ge0_a2 : c1995 ? jump_ge0_a2 : c1996 ? jump_ge0_a2 : ((c2055 || c2091) || c2090) ? jump_ge0_a2 : c1998 ? jump_ge0_a2 : c1999 ? jump_ge0_a2 : c2000 ? jump_ge0_a2 : c2001 ? jump_ge0_a2 : (c2199 || c2198) ? jump_ge0_a2 : (c2002 && !c927) ? jump_ge0_a2 : c1972 ? jump_ge0_a2 : 'bz; */
        /* jump_ge0_ip6 <= (c1971 && c889) ? jump_ge0_ip2 : ((c2004 || c2005) || c2006) ? jump_ge0_ip2 : c1974 ? jump_ge0_ip2 : c1975 ? jump_ge0_ip2 : c1976 ? jump_ge0_ip2 : c1977 ? jump_ge0_ip2 : c1978 ? jump_ge0_ip2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? jump_ge0_ip2 : (((c2019 || c2017) || c2018) || c2016) ? jump_ge0_ip2 : c1981 ? jump_ge0_ip2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? jump_ge0_ip5 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? jump_ge0_ip2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? jump_ge0_ip2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? jump_ge0_ip2 : (((c2038 || c2040) || c2037) || c2039) ? jump_ge0_ip2 : (c2041 || c2042) ? jump_ge0_ip2 : c1988 ? jump_ge0_ip2 : c1989 ? jump_ge0_ip2 : c1990 ? jump_ge0_ip2 : c1991 ? jump_ge0_ip2 : c1992 ? jump_ge0_ip2 : c1993 ? jump_ge0_ip2 : c1994 ? jump_ge0_ip2 : c1995 ? jump_ge0_ip2 : c1996 ? jump_ge0_ip2 : ((c2055 || c2091) || c2090) ? jump_ge0_ip2 : c1998 ? jump_ge0_ip2 : c1999 ? jump_ge0_ip2 : c2000 ? jump_ge0_ip2 : c2001 ? jump_ge0_ip2 : (c2199 || c2198) ? jump_ge0_ip2 : (c2002 && !c927) ? jump_ge0_ip2 : c1972 ? jump_ge0_ip2 : 'bz; */
        /* jump_ge0_phase9 <= (c1971 && c889) ? jump_ge0_phase2 : ((c2004 || c2005) || c2006) ? jump_ge0_phase2 : c1974 ? jump_ge0_phase2 : c1975 ? jump_ge0_phase2 : c1976 ? jump_ge0_phase2 : c1977 ? jump_ge0_phase2 : c1978 ? jump_ge0_phase2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? jump_ge0_phase2 : (((c2019 || c2017) || c2018) || c2016) ? jump_ge0_phase2 : c1981 ? jump_ge0_phase2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? jump_ge0_phase8 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? jump_ge0_phase2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? jump_ge0_phase2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? jump_ge0_phase2 : (((c2038 || c2040) || c2037) || c2039) ? jump_ge0_phase2 : (c2041 || c2042) ? jump_ge0_phase2 : c1988 ? jump_ge0_phase2 : c1989 ? jump_ge0_phase2 : c1990 ? jump_ge0_phase2 : c1991 ? jump_ge0_phase2 : c1992 ? jump_ge0_phase2 : c1993 ? jump_ge0_phase2 : c1994 ? jump_ge0_phase2 : c1995 ? jump_ge0_phase2 : c1996 ? jump_ge0_phase2 : ((c2055 || c2091) || c2090) ? jump_ge0_phase2 : c1998 ? jump_ge0_phase2 : c1999 ? jump_ge0_phase2 : c2000 ? jump_ge0_phase2 : c2001 ? jump_ge0_phase2 : (c2199 || c2198) ? jump_ge0_phase2 : (c2002 && !c927) ? jump_ge0_phase2 : c1972 ? jump_ge0_phase2 : 'bz; */
        /* jump_le0_a5 <= (c1971 && c889) ? jump_le0_a2 : ((c2004 || c2005) || c2006) ? jump_le0_a2 : c1974 ? jump_le0_a2 : c1975 ? jump_le0_a2 : c1976 ? jump_le0_a2 : c1977 ? jump_le0_a2 : c1978 ? jump_le0_a2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? jump_le0_a2 : (((c2019 || c2017) || c2018) || c2016) ? jump_le0_a2 : c1981 ? jump_le0_a2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? jump_le0_a2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? jump_le0_a4 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? jump_le0_a2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? jump_le0_a2 : (((c2038 || c2040) || c2037) || c2039) ? jump_le0_a2 : (c2041 || c2042) ? jump_le0_a2 : c1988 ? jump_le0_a2 : c1989 ? jump_le0_a2 : c1990 ? jump_le0_a2 : c1991 ? jump_le0_a2 : c1992 ? jump_le0_a2 : c1993 ? jump_le0_a2 : c1994 ? jump_le0_a2 : c1995 ? jump_le0_a2 : c1996 ? jump_le0_a2 : ((c2055 || c2091) || c2090) ? jump_le0_a2 : c1998 ? jump_le0_a2 : c1999 ? jump_le0_a2 : c2000 ? jump_le0_a2 : c2001 ? jump_le0_a2 : (c2199 || c2198) ? jump_le0_a2 : (c2002 && !c927) ? jump_le0_a2 : c1972 ? jump_le0_a2 : 'bz; */
        /* jump_le0_ip6 <= (c1971 && c889) ? jump_le0_ip2 : ((c2004 || c2005) || c2006) ? jump_le0_ip2 : c1974 ? jump_le0_ip2 : c1975 ? jump_le0_ip2 : c1976 ? jump_le0_ip2 : c1977 ? jump_le0_ip2 : c1978 ? jump_le0_ip2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? jump_le0_ip2 : (((c2019 || c2017) || c2018) || c2016) ? jump_le0_ip2 : c1981 ? jump_le0_ip2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? jump_le0_ip2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? jump_le0_ip5 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? jump_le0_ip2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? jump_le0_ip2 : (((c2038 || c2040) || c2037) || c2039) ? jump_le0_ip2 : (c2041 || c2042) ? jump_le0_ip2 : c1988 ? jump_le0_ip2 : c1989 ? jump_le0_ip2 : c1990 ? jump_le0_ip2 : c1991 ? jump_le0_ip2 : c1992 ? jump_le0_ip2 : c1993 ? jump_le0_ip2 : c1994 ? jump_le0_ip2 : c1995 ? jump_le0_ip2 : c1996 ? jump_le0_ip2 : ((c2055 || c2091) || c2090) ? jump_le0_ip2 : c1998 ? jump_le0_ip2 : c1999 ? jump_le0_ip2 : c2000 ? jump_le0_ip2 : c2001 ? jump_le0_ip2 : (c2199 || c2198) ? jump_le0_ip2 : (c2002 && !c927) ? jump_le0_ip2 : c1972 ? jump_le0_ip2 : 'bz; */
        /* jump_le0_phase9 <= (c1971 && c889) ? jump_le0_phase2 : ((c2004 || c2005) || c2006) ? jump_le0_phase2 : c1974 ? jump_le0_phase2 : c1975 ? jump_le0_phase2 : c1976 ? jump_le0_phase2 : c1977 ? jump_le0_phase2 : c1978 ? jump_le0_phase2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? jump_le0_phase2 : (((c2019 || c2017) || c2018) || c2016) ? jump_le0_phase2 : c1981 ? jump_le0_phase2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? jump_le0_phase2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? jump_le0_phase8 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? jump_le0_phase2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? jump_le0_phase2 : (((c2038 || c2040) || c2037) || c2039) ? jump_le0_phase2 : (c2041 || c2042) ? jump_le0_phase2 : c1988 ? jump_le0_phase2 : c1989 ? jump_le0_phase2 : c1990 ? jump_le0_phase2 : c1991 ? jump_le0_phase2 : c1992 ? jump_le0_phase2 : c1993 ? jump_le0_phase2 : c1994 ? jump_le0_phase2 : c1995 ? jump_le0_phase2 : c1996 ? jump_le0_phase2 : ((c2055 || c2091) || c2090) ? jump_le0_phase2 : c1998 ? jump_le0_phase2 : c1999 ? jump_le0_phase2 : c2000 ? jump_le0_phase2 : c2001 ? jump_le0_phase2 : (c2199 || c2198) ? jump_le0_phase2 : (c2002 && !c927) ? jump_le0_phase2 : c1972 ? jump_le0_phase2 : 'bz; */
        /* jump_ne0_a5 <= (c1971 && c889) ? jump_ne0_a2 : ((c2004 || c2005) || c2006) ? jump_ne0_a2 : c1974 ? jump_ne0_a2 : c1975 ? jump_ne0_a2 : c1976 ? jump_ne0_a2 : c1977 ? jump_ne0_a2 : c1978 ? jump_ne0_a2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? jump_ne0_a2 : (((c2019 || c2017) || c2018) || c2016) ? jump_ne0_a2 : c1981 ? jump_ne0_a2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? jump_ne0_a2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? jump_ne0_a2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? jump_ne0_a4 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? jump_ne0_a2 : (((c2038 || c2040) || c2037) || c2039) ? jump_ne0_a2 : (c2041 || c2042) ? jump_ne0_a2 : c1988 ? jump_ne0_a2 : c1989 ? jump_ne0_a2 : c1990 ? jump_ne0_a2 : c1991 ? jump_ne0_a2 : c1992 ? jump_ne0_a2 : c1993 ? jump_ne0_a2 : c1994 ? jump_ne0_a2 : c1995 ? jump_ne0_a2 : c1996 ? jump_ne0_a2 : ((c2055 || c2091) || c2090) ? jump_ne0_a2 : c1998 ? jump_ne0_a2 : c1999 ? jump_ne0_a2 : c2000 ? jump_ne0_a2 : c2001 ? jump_ne0_a2 : (c2199 || c2198) ? jump_ne0_a2 : (c2002 && !c927) ? jump_ne0_a2 : c1972 ? jump_ne0_a2 : 'bz; */
        /* jump_ne0_ip6 <= (c1971 && c889) ? jump_ne0_ip2 : ((c2004 || c2005) || c2006) ? jump_ne0_ip2 : c1974 ? jump_ne0_ip2 : c1975 ? jump_ne0_ip2 : c1976 ? jump_ne0_ip2 : c1977 ? jump_ne0_ip2 : c1978 ? jump_ne0_ip2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? jump_ne0_ip2 : (((c2019 || c2017) || c2018) || c2016) ? jump_ne0_ip2 : c1981 ? jump_ne0_ip2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? jump_ne0_ip2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? jump_ne0_ip2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? jump_ne0_ip5 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? jump_ne0_ip2 : (((c2038 || c2040) || c2037) || c2039) ? jump_ne0_ip2 : (c2041 || c2042) ? jump_ne0_ip2 : c1988 ? jump_ne0_ip2 : c1989 ? jump_ne0_ip2 : c1990 ? jump_ne0_ip2 : c1991 ? jump_ne0_ip2 : c1992 ? jump_ne0_ip2 : c1993 ? jump_ne0_ip2 : c1994 ? jump_ne0_ip2 : c1995 ? jump_ne0_ip2 : c1996 ? jump_ne0_ip2 : ((c2055 || c2091) || c2090) ? jump_ne0_ip2 : c1998 ? jump_ne0_ip2 : c1999 ? jump_ne0_ip2 : c2000 ? jump_ne0_ip2 : c2001 ? jump_ne0_ip2 : (c2199 || c2198) ? jump_ne0_ip2 : (c2002 && !c927) ? jump_ne0_ip2 : c1972 ? jump_ne0_ip2 : 'bz; */
        /* jump_ne0_phase9 <= (c1971 && c889) ? jump_ne0_phase2 : ((c2004 || c2005) || c2006) ? jump_ne0_phase2 : c1974 ? jump_ne0_phase2 : c1975 ? jump_ne0_phase2 : c1976 ? jump_ne0_phase2 : c1977 ? jump_ne0_phase2 : c1978 ? jump_ne0_phase2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? jump_ne0_phase2 : (((c2019 || c2017) || c2018) || c2016) ? jump_ne0_phase2 : c1981 ? jump_ne0_phase2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? jump_ne0_phase2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? jump_ne0_phase2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? jump_ne0_phase8 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? jump_ne0_phase2 : (((c2038 || c2040) || c2037) || c2039) ? jump_ne0_phase2 : (c2041 || c2042) ? jump_ne0_phase2 : c1988 ? jump_ne0_phase2 : c1989 ? jump_ne0_phase2 : c1990 ? jump_ne0_phase2 : c1991 ? jump_ne0_phase2 : c1992 ? jump_ne0_phase2 : c1993 ? jump_ne0_phase2 : c1994 ? jump_ne0_phase2 : c1995 ? jump_ne0_phase2 : c1996 ? jump_ne0_phase2 : ((c2055 || c2091) || c2090) ? jump_ne0_phase2 : c1998 ? jump_ne0_phase2 : c1999 ? jump_ne0_phase2 : c2000 ? jump_ne0_phase2 : c2001 ? jump_ne0_phase2 : (c2199 || c2198) ? jump_ne0_phase2 : (c2002 && !c927) ? jump_ne0_phase2 : c1972 ? jump_ne0_phase2 : 'bz; */
        /* lit0_ip5 <= (c1971 && c889) ? lit0_ip2 : ((c2004 || c2005) || c2006) ? lit0_ip4 : c1974 ? lit0_ip2 : c1975 ? lit0_ip2 : c1976 ? lit0_ip2 : c1977 ? lit0_ip2 : c1978 ? lit0_ip2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? lit0_ip2 : (((c2019 || c2017) || c2018) || c2016) ? lit0_ip2 : c1981 ? lit0_ip2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? lit0_ip2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? lit0_ip2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? lit0_ip2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? lit0_ip2 : (((c2038 || c2040) || c2037) || c2039) ? lit0_ip2 : (c2041 || c2042) ? lit0_ip2 : c1988 ? lit0_ip2 : c1989 ? lit0_ip2 : c1990 ? lit0_ip2 : c1991 ? lit0_ip2 : c1992 ? lit0_ip2 : c1993 ? lit0_ip2 : c1994 ? lit0_ip2 : c1995 ? lit0_ip2 : c1996 ? lit0_ip2 : ((c2055 || c2091) || c2090) ? lit0_ip2 : c1998 ? lit0_ip2 : c1999 ? lit0_ip2 : c2000 ? lit0_ip2 : c2001 ? lit0_ip2 : (c2199 || c2198) ? lit0_ip2 : (c2002 && !c927) ? lit0_ip2 : c1972 ? lit0_ip2 : 'bz; */
        /* lit0_phase7 <= (c1971 && c889) ? lit0_phase2 : ((c2004 || c2005) || c2006) ? lit0_phase6 : c1974 ? lit0_phase2 : c1975 ? lit0_phase2 : c1976 ? lit0_phase2 : c1977 ? lit0_phase2 : c1978 ? lit0_phase2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? lit0_phase2 : (((c2019 || c2017) || c2018) || c2016) ? lit0_phase2 : c1981 ? lit0_phase2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? lit0_phase2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? lit0_phase2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? lit0_phase2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? lit0_phase2 : (((c2038 || c2040) || c2037) || c2039) ? lit0_phase2 : (c2041 || c2042) ? lit0_phase2 : c1988 ? lit0_phase2 : c1989 ? lit0_phase2 : c1990 ? lit0_phase2 : c1991 ? lit0_phase2 : c1992 ? lit0_phase2 : c1993 ? lit0_phase2 : c1994 ? lit0_phase2 : c1995 ? lit0_phase2 : c1996 ? lit0_phase2 : ((c2055 || c2091) || c2090) ? lit0_phase2 : c1998 ? lit0_phase2 : c1999 ? lit0_phase2 : c2000 ? lit0_phase2 : c2001 ? lit0_phase2 : (c2199 || c2198) ? lit0_phase2 : (c2002 && !c927) ? lit0_phase2 : c1972 ? lit0_phase2 : 'bz; */
        /* loop0_ip6 <= (c1971 && c889) ? loop0_ip2 : ((c2004 || c2005) || c2006) ? loop0_ip2 : c1974 ? loop0_ip2 : c1975 ? loop0_ip2 : c1976 ? loop0_ip2 : c1977 ? loop0_ip2 : c1978 ? loop0_ip2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? loop0_ip5 : (((c2019 || c2017) || c2018) || c2016) ? loop0_ip2 : c1981 ? loop0_ip2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? loop0_ip2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? loop0_ip2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? loop0_ip2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? loop0_ip2 : (((c2038 || c2040) || c2037) || c2039) ? loop0_ip2 : (c2041 || c2042) ? loop0_ip2 : c1988 ? loop0_ip2 : c1989 ? loop0_ip2 : c1990 ? loop0_ip2 : c1991 ? loop0_ip2 : c1992 ? loop0_ip2 : c1993 ? loop0_ip2 : c1994 ? loop0_ip2 : c1995 ? loop0_ip2 : c1996 ? loop0_ip2 : ((c2055 || c2091) || c2090) ? loop0_ip2 : c1998 ? loop0_ip2 : c1999 ? loop0_ip2 : c2000 ? loop0_ip2 : c2001 ? loop0_ip2 : (c2199 || c2198) ? loop0_ip2 : (c2002 && !c927) ? loop0_ip2 : c1972 ? loop0_ip2 : 'bz; */
        /* loop0_phase9 <= (c1971 && c889) ? loop0_phase2 : ((c2004 || c2005) || c2006) ? loop0_phase2 : c1974 ? loop0_phase2 : c1975 ? loop0_phase2 : c1976 ? loop0_phase2 : c1977 ? loop0_phase2 : c1978 ? loop0_phase2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? loop0_phase8 : (((c2019 || c2017) || c2018) || c2016) ? loop0_phase2 : c1981 ? loop0_phase2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? loop0_phase2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? loop0_phase2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? loop0_phase2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? loop0_phase2 : (((c2038 || c2040) || c2037) || c2039) ? loop0_phase2 : (c2041 || c2042) ? loop0_phase2 : c1988 ? loop0_phase2 : c1989 ? loop0_phase2 : c1990 ? loop0_phase2 : c1991 ? loop0_phase2 : c1992 ? loop0_phase2 : c1993 ? loop0_phase2 : c1994 ? loop0_phase2 : c1995 ? loop0_phase2 : c1996 ? loop0_phase2 : ((c2055 || c2091) || c2090) ? loop0_phase2 : c1998 ? loop0_phase2 : c1999 ? loop0_phase2 : c2000 ? loop0_phase2 : c2001 ? loop0_phase2 : (c2199 || c2198) ? loop0_phase2 : (c2002 && !c927) ? loop0_phase2 : c1972 ? loop0_phase2 : 'bz; */
        /* point0_ip6 <= (c1971 && c889) ? point0_ip2 : ((c2004 || c2005) || c2006) ? point0_ip2 : c1974 ? point0_ip2 : c1975 ? point0_ip2 : c1976 ? point0_ip2 : c1977 ? point0_ip2 : c1978 ? point0_ip2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? point0_ip2 : (((c2019 || c2017) || c2018) || c2016) ? point0_ip2 : c1981 ? point0_ip2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? point0_ip2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? point0_ip2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? point0_ip2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? point0_ip2 : (((c2038 || c2040) || c2037) || c2039) ? point0_ip5 : (c2041 || c2042) ? point0_ip2 : c1988 ? point0_ip2 : c1989 ? point0_ip2 : c1990 ? point0_ip2 : c1991 ? point0_ip2 : c1992 ? point0_ip2 : c1993 ? point0_ip2 : c1994 ? point0_ip2 : c1995 ? point0_ip2 : c1996 ? point0_ip2 : ((c2055 || c2091) || c2090) ? point0_ip2 : c1998 ? point0_ip2 : c1999 ? point0_ip2 : c2000 ? point0_ip2 : c2001 ? point0_ip2 : (c2199 || c2198) ? point0_ip2 : (c2002 && !c927) ? point0_ip2 : c1972 ? point0_ip2 : 'bz; */
        /* point0_ip_saved5 <= (c1971 && c889) ? point0_ip_saved2 : ((c2004 || c2005) || c2006) ? point0_ip_saved2 : c1974 ? point0_ip_saved2 : c1975 ? point0_ip_saved2 : c1976 ? point0_ip_saved2 : c1977 ? point0_ip_saved2 : c1978 ? point0_ip_saved2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? point0_ip_saved2 : (((c2019 || c2017) || c2018) || c2016) ? point0_ip_saved2 : c1981 ? point0_ip_saved2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? point0_ip_saved2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? point0_ip_saved2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? point0_ip_saved2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? point0_ip_saved2 : (((c2038 || c2040) || c2037) || c2039) ? point0_ip_saved4 : (c2041 || c2042) ? point0_ip_saved2 : c1988 ? point0_ip_saved2 : c1989 ? point0_ip_saved2 : c1990 ? point0_ip_saved2 : c1991 ? point0_ip_saved2 : c1992 ? point0_ip_saved2 : c1993 ? point0_ip_saved2 : c1994 ? point0_ip_saved2 : c1995 ? point0_ip_saved2 : c1996 ? point0_ip_saved2 : ((c2055 || c2091) || c2090) ? point0_ip_saved2 : c1998 ? point0_ip_saved2 : c1999 ? point0_ip_saved2 : c2000 ? point0_ip_saved2 : c2001 ? point0_ip_saved2 : (c2199 || c2198) ? point0_ip_saved2 : (c2002 && !c927) ? point0_ip_saved2 : c1972 ? point0_ip_saved2 : 'bz; */
        /* point0_phase8 <= (c1971 && c889) ? point0_phase2 : ((c2004 || c2005) || c2006) ? point0_phase2 : c1974 ? point0_phase2 : c1975 ? point0_phase2 : c1976 ? point0_phase2 : c1977 ? point0_phase2 : c1978 ? point0_phase2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? point0_phase2 : (((c2019 || c2017) || c2018) || c2016) ? point0_phase2 : c1981 ? point0_phase2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? point0_phase2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? point0_phase2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? point0_phase2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? point0_phase2 : (((c2038 || c2040) || c2037) || c2039) ? point0_phase7 : (c2041 || c2042) ? point0_phase2 : c1988 ? point0_phase2 : c1989 ? point0_phase2 : c1990 ? point0_phase2 : c1991 ? point0_phase2 : c1992 ? point0_phase2 : c1993 ? point0_phase2 : c1994 ? point0_phase2 : c1995 ? point0_phase2 : c1996 ? point0_phase2 : ((c2055 || c2091) || c2090) ? point0_phase2 : c1998 ? point0_phase2 : c1999 ? point0_phase2 : c2000 ? point0_phase2 : c2001 ? point0_phase2 : (c2199 || c2198) ? point0_phase2 : (c2002 && !c927) ? point0_phase2 : c1972 ? point0_phase2 : 'bz; */
        /* stack0_pos43 <= (c1971 && c889) ? stack0_pos2 : ((c2004 || c2005) || c2006) ? stack0_pos4 : c1974 ? stack0_pos5 : c1975 ? stack0_pos6 : c1976 ? stack0_pos2 : c1977 ? stack0_pos7 : c1978 ? stack0_pos8 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? stack0_pos10 : (((c2019 || c2017) || c2018) || c2016) ? stack0_pos2 : c1981 ? stack0_pos2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? stack0_pos13 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? stack0_pos16 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? stack0_pos19 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? stack0_pos22 : (((c2038 || c2040) || c2037) || c2039) ? stack0_pos2 : (c2041 || c2042) ? stack0_pos25 : c1988 ? stack0_pos26 : c1989 ? stack0_pos27 : c1990 ? stack0_pos28 : c1991 ? stack0_pos2 : c1992 ? stack0_pos29 : c1993 ? stack0_pos30 : c1994 ? stack0_pos31 : c1995 ? stack0_pos32 : c1996 ? stack0_pos33 : ((c2055 || c2091) || c2090) ? stack0_pos35 : c1998 ? stack0_pos2 : c1999 ? stack0_pos2 : c2000 ? stack0_pos2 : c2001 ? stack0_pos37 : (c2199 || c2198) ? stack0_pos42 : (c2002 && !c927) ? stack0_pos2 : c1972 ? stack0_pos2 : 'bz; */
        /* stack0_second45 <= (c1971 && c889) ? stack0_second2 : ((c2004 || c2005) || c2006) ? stack0_second4 : c1974 ? stack0_top2 : c1975 ? stack0_second6 : c1976 ? stack0_top2 : c1977 ? stack0_second8 : c1978 ? stack0_top2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? stack0_second11 : (((c2019 || c2017) || c2018) || c2016) ? stack0_second2 : c1981 ? stack0_second2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? stack0_second14 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? stack0_second17 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? stack0_second20 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? stack0_second23 : (((c2038 || c2040) || c2037) || c2039) ? stack0_second2 : (c2041 || c2042) ? stack0_second26 : c1988 ? stack0_second27 : c1989 ? stack0_second28 : c1990 ? stack0_second29 : c1991 ? stack0_second30 : c1992 ? stack0_second31 : c1993 ? stack0_second32 : c1994 ? stack0_second33 : c1995 ? stack0_second34 : c1996 ? stack0_second35 : ((c2055 || c2091) || c2090) ? stack0_second37 : c1998 ? stack0_second2 : c1999 ? stack0_second2 : c2000 ? stack0_second2 : c2001 ? stack0_second39 : (c2199 || c2198) ? stack0_second44 : (c2002 && !c927) ? stack0_second2 : c1972 ? stack0_second2 : 'bz; */
        /* stack0_top59 <= (c1971 && c889) ? stack0_top2 : ((c2004 || c2005) || c2006) ? stack0_top4 : c1974 ? stack0_top2 : c1975 ? stack0_second2 : c1976 ? stack0_second2 : c1977 ? stack0_second2 : c1978 ? address0_top2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? stack0_top12 : (((c2019 || c2017) || c2018) || c2016) ? stack0_top2 : c1981 ? stack0_top2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? stack0_top15 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? stack0_top18 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? stack0_top21 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? stack0_top24 : (((c2038 || c2040) || c2037) || c2039) ? stack0_top26 : (c2041 || c2042) ? stack0_second2 : c1988 ? stack0_top31 : c1989 ? stack0_top33 : c1990 ? stack0_top35 : c1991 ? stack0_top36 : c1992 ? stack0_top38 : c1993 ? stack0_top40 : c1994 ? stack0_top42 : c1995 ? stack0_top44 : c1996 ? stack0_top46 : ((c2055 || c2091) || c2090) ? stack0_top48 : c1998 ? stack0_top49 : c1999 ? stack0_top50 : c2000 ? stack0_top51 : c2001 ? stack0_second38 : (c2199 || c2198) ? stack0_top58 : (c2002 && !c927) ? stack0_top2 : c1972 ? stack0_top2 : 'bz; */
        t11 <= (c1971 && c889) ? t11 : ((c2004 || c2005) || c2006) ? t11 : c1974 ? t11 : c1975 ? t11 : c1976 ? t11 : c1977 ? t11 : c1978 ? t11 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? t11 : (((c2019 || c2017) || c2018) || c2016) ? t11 : c1981 ? t11 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? t11 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? t11 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? t11 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? t11 : (((c2038 || c2040) || c2037) || c2039) ? t11 : (c2041 || c2042) ? t11 : c1988 ? stack0_top2 : c1989 ? stack0_top2 : c1990 ? stack0_top2 : c1991 ? t11 : c1992 ? stack0_top2 : c1993 ? stack0_top2 : c1994 ? stack0_top2 : c1995 ? stack0_top2 : c1996 ? stack0_top2 : ((c2055 || c2091) || c2090) ? t11 : c1998 ? t11 : c1999 ? t11 : c2000 ? stack0_top2 : c2001 ? t11 : (c2199 || c2198) ? t11 : (c2002 && !c927) ? t11 : c1972 ? t11 : 'bz;
        /* wr_flag4 <= (c1971 && c889) ? wr_flag2 : ((c2004 || c2005) || c2006) ? wr_flag2 : c1974 ? wr_flag2 : c1975 ? wr_flag2 : c1976 ? wr_flag2 : c1977 ? wr_flag2 : c1978 ? wr_flag2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? wr_flag2 : (((c2019 || c2017) || c2018) || c2016) ? wr_flag2 : c1981 ? wr_flag2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? wr_flag2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? wr_flag2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? wr_flag2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? wr_flag2 : (((c2038 || c2040) || c2037) || c2039) ? wr_flag2 : (c2041 || c2042) ? t2829 : c1988 ? wr_flag2 : c1989 ? wr_flag2 : c1990 ? wr_flag2 : c1991 ? wr_flag2 : c1992 ? wr_flag2 : c1993 ? wr_flag2 : c1994 ? wr_flag2 : c1995 ? wr_flag2 : c1996 ? wr_flag2 : ((c2055 || c2091) || c2090) ? wr_flag2 : c1998 ? wr_flag2 : c1999 ? wr_flag2 : c2000 ? wr_flag2 : c2001 ? wr_flag2 : (c2199 || c2198) ? wr_flag2 : (c2002 && !c927) ? wr_flag2 : c1972 ? wr_flag2 : 'bz; */
        /* wr_mem_addr4 <= (c1971 && c889) ? wr_mem_addr2 : ((c2004 || c2005) || c2006) ? wr_mem_addr2 : c1974 ? wr_mem_addr2 : c1975 ? wr_mem_addr2 : c1976 ? wr_mem_addr2 : c1977 ? wr_mem_addr2 : c1978 ? wr_mem_addr2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? wr_mem_addr2 : (((c2019 || c2017) || c2018) || c2016) ? wr_mem_addr2 : c1981 ? wr_mem_addr2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? wr_mem_addr2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? wr_mem_addr2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? wr_mem_addr2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? wr_mem_addr2 : (((c2038 || c2040) || c2037) || c2039) ? wr_mem_addr2 : (c2041 || c2042) ? t2830 : c1988 ? wr_mem_addr2 : c1989 ? wr_mem_addr2 : c1990 ? wr_mem_addr2 : c1991 ? wr_mem_addr2 : c1992 ? wr_mem_addr2 : c1993 ? wr_mem_addr2 : c1994 ? wr_mem_addr2 : c1995 ? wr_mem_addr2 : c1996 ? wr_mem_addr2 : ((c2055 || c2091) || c2090) ? wr_mem_addr2 : c1998 ? wr_mem_addr2 : c1999 ? wr_mem_addr2 : c2000 ? wr_mem_addr2 : c2001 ? wr_mem_addr2 : (c2199 || c2198) ? wr_mem_addr2 : (c2002 && !c927) ? wr_mem_addr2 : c1972 ? wr_mem_addr2 : 'bz; */
        /* wr_mem_data4 <= (c1971 && c889) ? wr_mem_data2 : ((c2004 || c2005) || c2006) ? wr_mem_data2 : c1974 ? wr_mem_data2 : c1975 ? wr_mem_data2 : c1976 ? wr_mem_data2 : c1977 ? wr_mem_data2 : c1978 ? wr_mem_data2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? wr_mem_data2 : (((c2019 || c2017) || c2018) || c2016) ? wr_mem_data2 : c1981 ? wr_mem_data2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? wr_mem_data2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? wr_mem_data2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? wr_mem_data2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? wr_mem_data2 : (((c2038 || c2040) || c2037) || c2039) ? wr_mem_data2 : (c2041 || c2042) ? t2831 : c1988 ? wr_mem_data2 : c1989 ? wr_mem_data2 : c1990 ? wr_mem_data2 : c1991 ? wr_mem_data2 : c1992 ? wr_mem_data2 : c1993 ? wr_mem_data2 : c1994 ? wr_mem_data2 : c1995 ? wr_mem_data2 : c1996 ? wr_mem_data2 : ((c2055 || c2091) || c2090) ? wr_mem_data2 : c1998 ? wr_mem_data2 : c1999 ? wr_mem_data2 : c2000 ? wr_mem_data2 : c2001 ? wr_mem_data2 : (c2199 || c2198) ? wr_mem_data2 : (c2002 && !c927) ? wr_mem_data2 : c1972 ? wr_mem_data2 : 'bz; */
        /* write_point0_addr5 <= (c1971 && c889) ? write_point0_addr2 : ((c2004 || c2005) || c2006) ? write_point0_addr2 : c1974 ? write_point0_addr2 : c1975 ? write_point0_addr2 : c1976 ? write_point0_addr2 : c1977 ? write_point0_addr2 : c1978 ? write_point0_addr2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? write_point0_addr2 : (((c2019 || c2017) || c2018) || c2016) ? write_point0_addr2 : c1981 ? write_point0_addr2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? write_point0_addr2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? write_point0_addr2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? write_point0_addr2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? write_point0_addr2 : (((c2038 || c2040) || c2037) || c2039) ? write_point0_addr2 : (c2041 || c2042) ? write_point0_addr4 : c1988 ? write_point0_addr2 : c1989 ? write_point0_addr2 : c1990 ? write_point0_addr2 : c1991 ? write_point0_addr2 : c1992 ? write_point0_addr2 : c1993 ? write_point0_addr2 : c1994 ? write_point0_addr2 : c1995 ? write_point0_addr2 : c1996 ? write_point0_addr2 : ((c2055 || c2091) || c2090) ? write_point0_addr2 : c1998 ? write_point0_addr2 : c1999 ? write_point0_addr2 : c2000 ? write_point0_addr2 : c2001 ? write_point0_addr2 : (c2199 || c2198) ? write_point0_addr2 : (c2002 && !c927) ? write_point0_addr2 : c1972 ? write_point0_addr2 : 'bz; */
        /* write_point0_data5 <= (c1971 && c889) ? write_point0_data2 : ((c2004 || c2005) || c2006) ? write_point0_data2 : c1974 ? write_point0_data2 : c1975 ? write_point0_data2 : c1976 ? write_point0_data2 : c1977 ? write_point0_data2 : c1978 ? write_point0_data2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? write_point0_data2 : (((c2019 || c2017) || c2018) || c2016) ? write_point0_data2 : c1981 ? write_point0_data2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? write_point0_data2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? write_point0_data2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? write_point0_data2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? write_point0_data2 : (((c2038 || c2040) || c2037) || c2039) ? write_point0_data2 : (c2041 || c2042) ? write_point0_data4 : c1988 ? write_point0_data2 : c1989 ? write_point0_data2 : c1990 ? write_point0_data2 : c1991 ? write_point0_data2 : c1992 ? write_point0_data2 : c1993 ? write_point0_data2 : c1994 ? write_point0_data2 : c1995 ? write_point0_data2 : c1996 ? write_point0_data2 : ((c2055 || c2091) || c2090) ? write_point0_data2 : c1998 ? write_point0_data2 : c1999 ? write_point0_data2 : c2000 ? write_point0_data2 : c2001 ? write_point0_data2 : (c2199 || c2198) ? write_point0_data2 : (c2002 && !c927) ? write_point0_data2 : c1972 ? write_point0_data2 : 'bz; */
        /* write_point0_ip5 <= (c1971 && c889) ? write_point0_ip2 : ((c2004 || c2005) || c2006) ? write_point0_ip2 : c1974 ? write_point0_ip2 : c1975 ? write_point0_ip2 : c1976 ? write_point0_ip2 : c1977 ? write_point0_ip2 : c1978 ? write_point0_ip2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? write_point0_ip2 : (((c2019 || c2017) || c2018) || c2016) ? write_point0_ip2 : c1981 ? write_point0_ip2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? write_point0_ip2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? write_point0_ip2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? write_point0_ip2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? write_point0_ip2 : (((c2038 || c2040) || c2037) || c2039) ? write_point0_ip2 : (c2041 || c2042) ? write_point0_ip4 : c1988 ? write_point0_ip2 : c1989 ? write_point0_ip2 : c1990 ? write_point0_ip2 : c1991 ? write_point0_ip2 : c1992 ? write_point0_ip2 : c1993 ? write_point0_ip2 : c1994 ? write_point0_ip2 : c1995 ? write_point0_ip2 : c1996 ? write_point0_ip2 : ((c2055 || c2091) || c2090) ? write_point0_ip2 : c1998 ? write_point0_ip2 : c1999 ? write_point0_ip2 : c2000 ? write_point0_ip2 : c2001 ? write_point0_ip2 : (c2199 || c2198) ? write_point0_ip2 : (c2002 && !c927) ? write_point0_ip2 : c1972 ? write_point0_ip2 : 'bz; */
        /* write_point0_phase6 <= (c1971 && c889) ? write_point0_phase2 : ((c2004 || c2005) || c2006) ? write_point0_phase2 : c1974 ? write_point0_phase2 : c1975 ? write_point0_phase2 : c1976 ? write_point0_phase2 : c1977 ? write_point0_phase2 : c1978 ? write_point0_phase2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? write_point0_phase2 : (((c2019 || c2017) || c2018) || c2016) ? write_point0_phase2 : c1981 ? write_point0_phase2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? write_point0_phase2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? write_point0_phase2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? write_point0_phase2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? write_point0_phase2 : (((c2038 || c2040) || c2037) || c2039) ? write_point0_phase2 : (c2041 || c2042) ? write_point0_phase5 : c1988 ? write_point0_phase2 : c1989 ? write_point0_phase2 : c1990 ? write_point0_phase2 : c1991 ? write_point0_phase2 : c1992 ? write_point0_phase2 : c1993 ? write_point0_phase2 : c1994 ? write_point0_phase2 : c1995 ? write_point0_phase2 : c1996 ? write_point0_phase2 : ((c2055 || c2091) || c2090) ? write_point0_phase2 : c1998 ? write_point0_phase2 : c1999 ? write_point0_phase2 : c2000 ? write_point0_phase2 : c2001 ? write_point0_phase2 : (c2199 || c2198) ? write_point0_phase2 : (c2002 && !c927) ? write_point0_phase2 : c1972 ? write_point0_phase2 : 'bz; */
        /* zero_pop_return0_ip6 <= (c1971 && c889) ? zero_pop_return0_ip2 : ((c2004 || c2005) || c2006) ? zero_pop_return0_ip2 : c1974 ? zero_pop_return0_ip2 : c1975 ? zero_pop_return0_ip2 : c1976 ? zero_pop_return0_ip2 : c1977 ? zero_pop_return0_ip2 : c1978 ? zero_pop_return0_ip2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? zero_pop_return0_ip2 : (((c2019 || c2017) || c2018) || c2016) ? zero_pop_return0_ip2 : c1981 ? zero_pop_return0_ip2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? zero_pop_return0_ip2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? zero_pop_return0_ip2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? zero_pop_return0_ip2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? zero_pop_return0_ip2 : (((c2038 || c2040) || c2037) || c2039) ? zero_pop_return0_ip2 : (c2041 || c2042) ? zero_pop_return0_ip2 : c1988 ? zero_pop_return0_ip2 : c1989 ? zero_pop_return0_ip2 : c1990 ? zero_pop_return0_ip2 : c1991 ? zero_pop_return0_ip2 : c1992 ? zero_pop_return0_ip2 : c1993 ? zero_pop_return0_ip2 : c1994 ? zero_pop_return0_ip2 : c1995 ? zero_pop_return0_ip2 : c1996 ? zero_pop_return0_ip2 : ((c2055 || c2091) || c2090) ? zero_pop_return0_ip5 : c1998 ? zero_pop_return0_ip2 : c1999 ? zero_pop_return0_ip2 : c2000 ? zero_pop_return0_ip2 : c2001 ? zero_pop_return0_ip2 : (c2199 || c2198) ? zero_pop_return0_ip2 : (c2002 && !c927) ? zero_pop_return0_ip2 : c1972 ? zero_pop_return0_ip2 : 'bz; */
        /* zero_pop_return0_phase6 <= (c1971 && c889) ? zero_pop_return0_phase2 : ((c2004 || c2005) || c2006) ? zero_pop_return0_phase2 : c1974 ? zero_pop_return0_phase2 : c1975 ? zero_pop_return0_phase2 : c1976 ? zero_pop_return0_phase2 : c1977 ? zero_pop_return0_phase2 : c1978 ? zero_pop_return0_phase2 : ((((c2013 || c2015) || c2014) || c2124) || c2125) ? zero_pop_return0_phase2 : (((c2019 || c2017) || c2018) || c2016) ? zero_pop_return0_phase2 : c1981 ? zero_pop_return0_phase2 : ((((c2023 || c2024) || c2021) || c2126) || c2127) ? zero_pop_return0_phase2 : ((((c2028 || c2027) || c2025) || c2128) || c2129) ? zero_pop_return0_phase2 : ((((c2031 || c2032) || c2029) || c2130) || c2131) ? zero_pop_return0_phase2 : ((((c2036 || c2035) || c2033) || c2132) || c2133) ? zero_pop_return0_phase2 : (((c2038 || c2040) || c2037) || c2039) ? zero_pop_return0_phase2 : (c2041 || c2042) ? zero_pop_return0_phase2 : c1988 ? zero_pop_return0_phase2 : c1989 ? zero_pop_return0_phase2 : c1990 ? zero_pop_return0_phase2 : c1991 ? zero_pop_return0_phase2 : c1992 ? zero_pop_return0_phase2 : c1993 ? zero_pop_return0_phase2 : c1994 ? zero_pop_return0_phase2 : c1995 ? zero_pop_return0_phase2 : c1996 ? zero_pop_return0_phase2 : ((c2055 || c2091) || c2090) ? zero_pop_return0_phase5 : c1998 ? zero_pop_return0_phase2 : c1999 ? zero_pop_return0_phase2 : c2000 ? zero_pop_return0_phase2 : c2001 ? zero_pop_return0_phase2 : (c2199 || c2198) ? zero_pop_return0_phase2 : (c2002 && !c927) ? zero_pop_return0_phase2 : c1972 ? zero_pop_return0_phase2 : 'bz; */
        /* c920 <= (wr_flag4 != 0); */
        /* c2200 <= (c886 && c920); */
        retro_main_state <= retro_main_L1_b178_S1;
      end
      retro_main_L1_b178_S1: begin
        if (c920) begin
          memory_addr <= wr_mem_addr4;
          memory_we <= 1;
          memory_req <= 1;
          memory_d <= wr_mem_data4;
          /* c3450 <= (c886 && c920); */
          retro_main_state <= retro_main_L1_ifthen179_S1;
        end else begin
          opcode2 <= opcode4;
          /* c921 <= (done_flag13 != 0); */
          address0_pos2 <= address0_pos9;
          address0_second2 <= address0_second9;
          address0_top2 <= address0_top9;
          done_flag2 <= done_flag13;
          jump0_ip2 <= jump0_ip6;
          jump0_phase2 <= jump0_phase8;
          jump_eq0_a2 <= jump_eq0_a5;
          jump_eq0_ip2 <= jump_eq0_ip6;
          jump_eq0_phase2 <= jump_eq0_phase9;
          jump_ge0_a2 <= jump_ge0_a5;
          jump_ge0_ip2 <= jump_ge0_ip6;
          jump_ge0_phase2 <= jump_ge0_phase9;
          jump_le0_a2 <= jump_le0_a5;
          jump_le0_ip2 <= jump_le0_ip6;
          jump_le0_phase2 <= jump_le0_phase9;
          jump_ne0_a2 <= jump_ne0_a5;
          jump_ne0_ip2 <= jump_ne0_ip6;
          jump_ne0_phase2 <= jump_ne0_phase9;
          lit0_ip2 <= lit0_ip5;
          lit0_phase2 <= lit0_phase7;
          loop0_ip2 <= loop0_ip6;
          loop0_phase2 <= loop0_phase9;
          point0_ip2 <= point0_ip6;
          point0_ip_saved2 <= point0_ip_saved5;
          point0_phase2 <= point0_phase8;
          stack0_pos2 <= stack0_pos43;
          stack0_second2 <= stack0_second45;
          stack0_top2 <= stack0_top59;
          wr_mem_addr2 <= wr_mem_addr4;
          wr_mem_data2 <= wr_mem_data4;
          write_point0_addr2 <= write_point0_addr5;
          write_point0_data2 <= write_point0_data5;
          write_point0_ip2 <= write_point0_ip5;
          write_point0_phase2 <= write_point0_phase6;
          zero_pop_return0_ip2 <= zero_pop_return0_ip6;
          zero_pop_return0_phase2 <= zero_pop_return0_phase6;
          /* c2201 <= (c886 && c921); */
          /* wr_flag6 <= c2200 ? 0 : (c886 && !c920) ? wr_flag4 : 'bz; */
          wr_flag2 <= wr_flag6;
          retro_main_state <= retro_main_L1_b183_S1;
        end
      end
      retro_main_L1_ifthen179_S1: begin
        memory_req <= 0;
        retro_main_state <= retro_main_L1_b183_S0;
      end
      retro_main_L1_b183_S0: begin
        opcode2 <= opcode4;
        /* c921 <= (done_flag13 != 0); */
        address0_pos2 <= address0_pos9;
        address0_second2 <= address0_second9;
        address0_top2 <= address0_top9;
        done_flag2 <= done_flag13;
        jump0_ip2 <= jump0_ip6;
        jump0_phase2 <= jump0_phase8;
        jump_eq0_a2 <= jump_eq0_a5;
        jump_eq0_ip2 <= jump_eq0_ip6;
        jump_eq0_phase2 <= jump_eq0_phase9;
        jump_ge0_a2 <= jump_ge0_a5;
        jump_ge0_ip2 <= jump_ge0_ip6;
        jump_ge0_phase2 <= jump_ge0_phase9;
        jump_le0_a2 <= jump_le0_a5;
        jump_le0_ip2 <= jump_le0_ip6;
        jump_le0_phase2 <= jump_le0_phase9;
        jump_ne0_a2 <= jump_ne0_a5;
        jump_ne0_ip2 <= jump_ne0_ip6;
        jump_ne0_phase2 <= jump_ne0_phase9;
        lit0_ip2 <= lit0_ip5;
        lit0_phase2 <= lit0_phase7;
        loop0_ip2 <= loop0_ip6;
        loop0_phase2 <= loop0_phase9;
        point0_ip2 <= point0_ip6;
        point0_ip_saved2 <= point0_ip_saved5;
        point0_phase2 <= point0_phase8;
        stack0_pos2 <= stack0_pos43;
        stack0_second2 <= stack0_second45;
        stack0_top2 <= stack0_top59;
        wr_mem_addr2 <= wr_mem_addr4;
        wr_mem_data2 <= wr_mem_data4;
        write_point0_addr2 <= write_point0_addr5;
        write_point0_data2 <= write_point0_data5;
        write_point0_ip2 <= write_point0_ip5;
        write_point0_phase2 <= write_point0_phase6;
        zero_pop_return0_ip2 <= zero_pop_return0_ip6;
        zero_pop_return0_phase2 <= zero_pop_return0_phase6;
        /* c2201 <= (c886 && c921); */
        /* wr_flag6 <= c2200 ? 0 : (c886 && !c920) ? wr_flag4 : 'bz; */
        wr_flag2 <= wr_flag6;
        retro_main_state <= retro_main_L1_b183_S1;
      end
      retro_main_L1_b183_S1: begin
        /* ip17 <= (ip16 + 1); */
        /* ip18 <= c2201 ? ip17 : (c886 && !c921) ? ip16 : 'bz; */
        ip2 <= ip18;
        retro_main_state <= retro_main_L1_while2_S0;
      end
      endcase
    end
  end
  

endmodule

