module retro_main
  (
    input wire clk,
    input wire rst,
    input wire retro_main_ready,
    input wire retro_main_accept,
    output reg retro_main_valid,
    input wire signed [31:0] retro_main_in_memory_q,
    input wire [14:0] retro_main_in_memory_len,
    output wire signed [14:0] retro_main_in_memory_addr,
    output wire signed [31:0] retro_main_in_memory_d,
    output wire retro_main_in_memory_we,
    output wire retro_main_in_memory_req,
    input wire signed [31:0] retro_main_in_io_ports_q,
    input wire [4:0] retro_main_in_io_ports_len,
    output wire signed [4:0] retro_main_in_io_ports_addr,
    output wire signed [31:0] retro_main_in_io_ports_d,
    output wire retro_main_in_io_ports_we,
    output wire retro_main_in_io_ports_req
  );

  //localparams
  localparam retro_main_b1_INIT = 0;
  localparam retro_main_b1_S0 = 1;
  localparam retro_main_b1_S1 = 2;
  localparam retro_main_b1_S2 = 3;
  localparam retro_main_b1_S3 = 4;
  localparam retro_main_b1_S4 = 5;
  localparam retro_main_b1_S5 = 6;
  localparam retro_main_b1_S6 = 7;
  localparam retro_main_b1_S7 = 8;
  localparam retro_main_b1_S8 = 9;
  localparam retro_main_b1_S9 = 10;
  localparam retro_main_b1_S10 = 11;
  localparam retro_main_b1_S11 = 12;
  localparam retro_main_b1_S12 = 13;
  localparam retro_main_b1_S13 = 14;
  localparam retro_main_b1_S14 = 15;
  localparam retro_main_b1_S15 = 16;
  localparam retro_main_b1_S16 = 17;
  localparam retro_main_b1_S17 = 18;
  localparam retro_main_b1_S18 = 19;
  localparam retro_main_b1_S19 = 20;
  localparam retro_main_b1_S20 = 21;
  localparam retro_main_b1_S21 = 22;
  localparam retro_main_b1_S22 = 23;
  localparam retro_main_b1_S23 = 24;
  localparam retro_main_b1_S24 = 25;
  localparam retro_main_b1_S25 = 26;
  localparam retro_main_b1_S26 = 27;
  localparam retro_main_b1_S27 = 28;
  localparam retro_main_b1_S28 = 29;
  localparam retro_main_b1_S29 = 30;
  localparam retro_main_b1_S30 = 31;
  localparam retro_main_b1_S31 = 32;
  localparam retro_main_b1_S32 = 33;
  localparam retro_main_b1_S33 = 34;
  localparam retro_main_b1_S34 = 35;
  localparam retro_main_b1_S35 = 36;
  localparam retro_main_b1_S36 = 37;
  localparam retro_main_b1_S37 = 38;
  localparam retro_main_b1_S38 = 39;
  localparam retro_main_b1_S39 = 40;
  localparam retro_main_b1_S40 = 41;
  localparam retro_main_b1_S41 = 42;
  localparam retro_main_b1_S42 = 43;
  localparam retro_main_b1_S43 = 44;
  localparam retro_main_b1_S44 = 45;
  localparam retro_main_b1_S45 = 46;
  localparam retro_main_b1_S46 = 47;
  localparam retro_main_b1_S47 = 48;
  localparam retro_main_b1_S48 = 49;
  localparam retro_main_b1_S49 = 50;
  localparam retro_main_b1_S50 = 51;
  localparam retro_main_b1_S51 = 52;
  localparam retro_main_b1_S52 = 53;
  localparam retro_main_b1_S53 = 54;
  localparam retro_main_b1_S54 = 55;
  localparam retro_main_b1_S55 = 56;
  localparam retro_main_b1_S56 = 57;
  localparam retro_main_b1_S57 = 58;
  localparam retro_main_b1_S58 = 59;
  localparam retro_main_b1_S59 = 60;
  localparam retro_main_b1_S60 = 61;
  localparam retro_main_b1_S61 = 62;
  localparam retro_main_b1_S62 = 63;
  localparam retro_main_b1_S63 = 64;
  localparam retro_main_b1_S64 = 65;
  localparam retro_main_b1_S65 = 66;
  localparam retro_main_b1_S66 = 67;
  localparam retro_main_b1_S67 = 68;
  localparam retro_main_b1_S68 = 69;
  localparam retro_main_b1_S69 = 70;
  localparam retro_main_b1_S70 = 71;
  localparam retro_main_b1_S71 = 72;
  localparam retro_main_b1_S72 = 73;
  localparam retro_main_b1_S73 = 74;
  localparam retro_main_b1_S74 = 75;
  localparam retro_main_b1_S75 = 76;
  localparam retro_main_b1_S76 = 77;
  localparam retro_main_b1_S77 = 78;
  localparam retro_main_b1_S78 = 79;
  localparam retro_main_b1_S79 = 80;
  localparam retro_main_b1_S80 = 81;
  localparam retro_main_b1_S81 = 82;
  localparam retro_main_b1_S82 = 83;
  localparam retro_main_b1_S83 = 84;
  localparam retro_main_b1_S84 = 85;
  localparam retro_main_b1_S85 = 86;
  localparam retro_main_b1_S86 = 87;
  localparam retro_main_b1_S87 = 88;
  localparam retro_main_b1_S88 = 89;
  localparam retro_main_b1_S89 = 90;
  localparam retro_main_b1_S90 = 91;
  localparam retro_main_b1_S91 = 92;
  localparam retro_main_b1_S92 = 93;
  localparam retro_main_b1_S93 = 94;
  localparam retro_main_b1_S94 = 95;
  localparam retro_main_b1_S95 = 96;
  localparam retro_main_b1_S96 = 97;
  localparam retro_main_b1_S97 = 98;
  localparam retro_main_b1_S98 = 99;
  localparam retro_main_b1_S99 = 100;
  localparam retro_main_b1_S100 = 101;
  localparam retro_main_b1_S101 = 102;
  localparam retro_main_b1_S102 = 103;
  localparam retro_main_b1_S103 = 104;
  localparam retro_main_b1_S104 = 105;
  localparam retro_main_b1_S105 = 106;
  localparam retro_main_b1_S106 = 107;
  localparam retro_main_b1_S107 = 108;
  localparam retro_main_b1_S108 = 109;
  localparam retro_main_b1_S109 = 110;
  localparam retro_main_b1_S110 = 111;
  localparam retro_main_b1_S111 = 112;
  localparam retro_main_b1_S112 = 113;
  localparam retro_main_b1_S113 = 114;
  localparam retro_main_b1_S114 = 115;
  localparam retro_main_b1_S115 = 116;
  localparam retro_main_b1_S116 = 117;
  localparam retro_main_b1_S117 = 118;
  localparam retro_main_b1_S118 = 119;
  localparam retro_main_b1_S119 = 120;
  localparam retro_main_b1_S120 = 121;
  localparam retro_main_b1_S121 = 122;
  localparam retro_main_b1_S122 = 123;
  localparam retro_main_b1_S123 = 124;
  localparam retro_main_b1_S124 = 125;
  localparam retro_main_b1_S125 = 126;
  localparam retro_main_b1_S126 = 127;
  localparam retro_main_b1_S127 = 128;
  localparam retro_main_b1_S128 = 129;
  localparam retro_main_b1_S129 = 130;
  localparam retro_main_b1_S130 = 131;
  localparam retro_main_b1_S131 = 132;
  localparam retro_main_b1_S132 = 133;
  localparam retro_main_b1_S133 = 134;
  localparam retro_main_b1_S134 = 135;
  localparam retro_main_b1_S135 = 136;
  localparam retro_main_b1_S136 = 137;
  localparam retro_main_b1_S137 = 138;
  localparam retro_main_b1_S138 = 139;
  localparam retro_main_b1_S139 = 140;
  localparam retro_main_b1_S140 = 141;
  localparam retro_main_b1_S141 = 142;
  localparam retro_main_b1_S142 = 143;
  localparam retro_main_b1_S143 = 144;
  localparam retro_main_b1_S144 = 145;
  localparam retro_main_b1_S145 = 146;
  localparam retro_main_b1_S146 = 147;
  localparam retro_main_b1_S147 = 148;
  localparam retro_main_b1_S148 = 149;
  localparam retro_main_b1_S149 = 150;
  localparam retro_main_b1_S150 = 151;
  localparam retro_main_b1_S151 = 152;
  localparam retro_main_b1_S152 = 153;
  localparam retro_main_b1_S153 = 154;
  localparam retro_main_b1_S154 = 155;
  localparam retro_main_b1_S155 = 156;
  localparam retro_main_b1_S156 = 157;
  localparam retro_main_b1_S157 = 158;
  localparam retro_main_b1_S158 = 159;
  localparam retro_main_b1_S159 = 160;
  localparam retro_main_b1_S160 = 161;
  localparam retro_main_b1_S161 = 162;
  localparam retro_main_b1_S162 = 163;
  localparam retro_main_b1_S163 = 164;
  localparam retro_main_b1_S164 = 165;
  localparam retro_main_b1_S165 = 166;
  localparam retro_main_b1_S166 = 167;
  localparam retro_main_b1_S167 = 168;
  localparam retro_main_b1_S168 = 169;
  localparam retro_main_b1_S169 = 170;
  localparam retro_main_b1_S170 = 171;
  localparam retro_main_b1_S171 = 172;
  localparam retro_main_b1_S172 = 173;
  localparam retro_main_b1_S173 = 174;
  localparam retro_main_b1_S174 = 175;
  localparam retro_main_b1_S175 = 176;
  localparam retro_main_b1_S176 = 177;
  localparam retro_main_b1_S177 = 178;
  localparam retro_main_b1_S178 = 179;
  localparam retro_main_b1_S179 = 180;
  localparam retro_main_b1_S180 = 181;
  localparam retro_main_b1_S181 = 182;
  localparam retro_main_b1_S182 = 183;
  localparam retro_main_b1_S183 = 184;
  localparam retro_main_b1_S184 = 185;
  localparam retro_main_b1_S185 = 186;
  localparam retro_main_b1_S186 = 187;
  localparam retro_main_b1_S187 = 188;
  localparam retro_main_b1_S188 = 189;
  localparam retro_main_b1_S189 = 190;
  localparam retro_main_b1_S190 = 191;
  localparam retro_main_b1_S191 = 192;
  localparam retro_main_b1_S192 = 193;
  localparam retro_main_b1_S193 = 194;
  localparam retro_main_b1_S194 = 195;
  localparam retro_main_b1_S195 = 196;
  localparam retro_main_b1_S196 = 197;
  localparam retro_main_b1_S197 = 198;
  localparam retro_main_b1_S198 = 199;
  localparam retro_main_b1_S199 = 200;
  localparam retro_main_b1_S200 = 201;
  localparam retro_main_b1_S201 = 202;
  localparam retro_main_b1_S202 = 203;
  localparam retro_main_b1_S203 = 204;
  localparam retro_main_b1_S204 = 205;
  localparam retro_main_b1_S205 = 206;
  localparam retro_main_b1_S206 = 207;
  localparam retro_main_b1_S207 = 208;
  localparam retro_main_b1_S208 = 209;
  localparam retro_main_b1_S209 = 210;
  localparam retro_main_b1_S210 = 211;
  localparam retro_main_b1_S211 = 212;
  localparam retro_main_b1_S212 = 213;
  localparam retro_main_b1_S213 = 214;
  localparam retro_main_b1_S214 = 215;
  localparam retro_main_b1_S215 = 216;
  localparam retro_main_b1_S216 = 217;
  localparam retro_main_b1_S217 = 218;
  localparam retro_main_b1_S218 = 219;
  localparam retro_main_b1_S219 = 220;
  localparam retro_main_b1_S220 = 221;
  localparam retro_main_b1_S221 = 222;
  localparam retro_main_b1_S222 = 223;
  localparam retro_main_b1_S223 = 224;
  localparam retro_main_b1_S224 = 225;
  localparam retro_main_b1_S225 = 226;
  localparam retro_main_b1_S226 = 227;
  localparam retro_main_b1_S227 = 228;
  localparam retro_main_b1_S228 = 229;
  localparam retro_main_b1_S229 = 230;
  localparam retro_main_b1_S230 = 231;
  localparam retro_main_b1_S231 = 232;
  localparam retro_main_b1_S232 = 233;
  localparam retro_main_b1_S233 = 234;
  localparam retro_main_b1_S234 = 235;
  localparam retro_main_b1_S235 = 236;
  localparam retro_main_b1_S236 = 237;
  localparam retro_main_b1_S237 = 238;
  localparam retro_main_b1_S238 = 239;
  localparam retro_main_b1_S239 = 240;
  localparam retro_main_b1_S240 = 241;
  localparam retro_main_b1_S241 = 242;
  localparam retro_main_b1_S242 = 243;
  localparam retro_main_b1_S243 = 244;
  localparam retro_main_b1_S244 = 245;
  localparam retro_main_b1_S245 = 246;
  localparam retro_main_b1_S246 = 247;
  localparam retro_main_b1_S247 = 248;
  localparam retro_main_b1_S248 = 249;
  localparam retro_main_b1_S249 = 250;
  localparam retro_main_b1_S250 = 251;
  localparam retro_main_b1_S251 = 252;
  localparam retro_main_b1_S252 = 253;
  localparam retro_main_b1_S253 = 254;
  localparam retro_main_b1_S254 = 255;
  localparam retro_main_b1_S255 = 256;
  localparam retro_main_b1_S256 = 257;
  localparam retro_main_b1_S257 = 258;
  localparam retro_main_b1_S258 = 259;
  localparam retro_main_b1_S259 = 260;
  localparam retro_main_b1_S260 = 261;
  localparam retro_main_b1_S261 = 262;
  localparam retro_main_b1_S262 = 263;
  localparam retro_main_b1_S263 = 264;
  localparam retro_main_b1_S264 = 265;
  localparam retro_main_b1_S265 = 266;
  localparam retro_main_b1_S266 = 267;
  localparam retro_main_b1_S267 = 268;
  localparam retro_main_b1_S268 = 269;
  localparam retro_main_b1_S269 = 270;
  localparam retro_main_b1_S270 = 271;
  localparam retro_main_b1_S271 = 272;
  localparam retro_main_b1_S272 = 273;
  localparam retro_main_b1_S273 = 274;
  localparam retro_main_b1_S274 = 275;
  localparam retro_main_b1_S275 = 276;
  localparam retro_main_b1_S276 = 277;
  localparam retro_main_b1_S277 = 278;
  localparam retro_main_b1_S278 = 279;
  localparam retro_main_b1_S279 = 280;
  localparam retro_main_b1_S280 = 281;
  localparam retro_main_b1_S281 = 282;
  localparam retro_main_b1_S282 = 283;
  localparam retro_main_b1_S283 = 284;
  localparam retro_main_b1_S284 = 285;
  localparam retro_main_b1_S285 = 286;
  localparam retro_main_b1_S286 = 287;
  localparam retro_main_b1_S287 = 288;
  localparam retro_main_b1_S288 = 289;
  localparam retro_main_b1_S289 = 290;
  localparam retro_main_b1_S290 = 291;
  localparam retro_main_b1_S291 = 292;
  localparam retro_main_b1_S292 = 293;
  localparam retro_main_b1_S293 = 294;
  localparam retro_main_b1_S294 = 295;
  localparam retro_main_b1_S295 = 296;
  localparam retro_main_b1_S296 = 297;
  localparam retro_main_b1_S297 = 298;
  localparam retro_main_b1_S298 = 299;
  localparam retro_main_b1_S299 = 300;
  localparam retro_main_b1_S300 = 301;
  localparam retro_main_b1_S301 = 302;
  localparam retro_main_b1_S302 = 303;
  localparam retro_main_b1_S303 = 304;
  localparam retro_main_b1_S304 = 305;
  localparam retro_main_b1_S305 = 306;
  localparam retro_main_b1_S306 = 307;
  localparam retro_main_b1_S307 = 308;
  localparam retro_main_b1_S308 = 309;
  localparam retro_main_b1_S309 = 310;
  localparam retro_main_b1_S310 = 311;
  localparam retro_main_b1_S311 = 312;
  localparam retro_main_b1_S312 = 313;
  localparam retro_main_b1_S313 = 314;
  localparam retro_main_b1_S314 = 315;
  localparam retro_main_b1_S315 = 316;
  localparam retro_main_b1_S316 = 317;
  localparam retro_main_b1_S317 = 318;
  localparam retro_main_b1_S318 = 319;
  localparam retro_main_b1_S319 = 320;
  localparam retro_main_b1_S320 = 321;
  localparam retro_main_b1_S321 = 322;
  localparam retro_main_b1_S322 = 323;
  localparam retro_main_b1_S323 = 324;
  localparam retro_main_b1_S324 = 325;
  localparam retro_main_b1_S325 = 326;
  localparam retro_main_b1_S326 = 327;
  localparam retro_main_b1_S327 = 328;
  localparam retro_main_b1_S328 = 329;
  localparam retro_main_b1_S329 = 330;
  localparam retro_main_b1_S330 = 331;
  localparam retro_main_b1_S331 = 332;
  localparam retro_main_b1_S332 = 333;
  localparam retro_main_b1_S333 = 334;
  localparam retro_main_b1_S334 = 335;
  localparam retro_main_b1_S335 = 336;
  localparam retro_main_b1_S336 = 337;
  localparam retro_main_b1_S337 = 338;
  localparam retro_main_b1_S338 = 339;
  localparam retro_main_b1_S339 = 340;
  localparam retro_main_b1_S340 = 341;
  localparam retro_main_b1_S341 = 342;
  localparam retro_main_b1_S342 = 343;
  localparam retro_main_b1_S343 = 344;
  localparam retro_main_b1_S344 = 345;
  localparam retro_main_b1_S345 = 346;
  localparam retro_main_b1_S346 = 347;
  localparam retro_main_b1_S347 = 348;
  localparam retro_main_b1_S348 = 349;
  localparam retro_main_b1_S349 = 350;
  localparam retro_main_b1_S350 = 351;
  localparam retro_main_b1_S351 = 352;
  localparam retro_main_b1_S352 = 353;
  localparam retro_main_b1_S353 = 354;
  localparam retro_main_b1_S354 = 355;
  localparam retro_main_b1_S355 = 356;
  localparam retro_main_b1_S356 = 357;
  localparam retro_main_b1_S357 = 358;
  localparam retro_main_b1_S358 = 359;
  localparam retro_main_b1_S359 = 360;
  localparam retro_main_b1_S360 = 361;
  localparam retro_main_b1_S361 = 362;
  localparam retro_main_b1_S362 = 363;
  localparam retro_main_b1_S363 = 364;
  localparam retro_main_b1_S364 = 365;
  localparam retro_main_b1_S365 = 366;
  localparam retro_main_b1_S366 = 367;
  localparam retro_main_b1_S367 = 368;
  localparam retro_main_b1_S368 = 369;
  localparam retro_main_b1_S369 = 370;
  localparam retro_main_b1_S370 = 371;
  localparam retro_main_b1_S371 = 372;
  localparam retro_main_b1_S372 = 373;
  localparam retro_main_b1_S373 = 374;
  localparam retro_main_b1_S374 = 375;
  localparam retro_main_b1_S375 = 376;
  localparam retro_main_b1_S376 = 377;
  localparam retro_main_b1_S377 = 378;
  localparam retro_main_b1_S378 = 379;
  localparam retro_main_b1_S379 = 380;
  localparam retro_main_b1_S380 = 381;
  localparam retro_main_b1_S381 = 382;
  localparam retro_main_b1_S382 = 383;
  localparam retro_main_b1_S383 = 384;
  localparam retro_main_b1_S384 = 385;
  localparam retro_main_b1_S385 = 386;
  localparam retro_main_b1_S386 = 387;
  localparam retro_main_b1_S387 = 388;
  localparam retro_main_b1_S388 = 389;
  localparam retro_main_b1_S389 = 390;
  localparam retro_main_b1_S390 = 391;
  localparam retro_main_b1_S391 = 392;
  localparam retro_main_b1_S392 = 393;
  localparam retro_main_b1_S393 = 394;
  localparam retro_main_b1_S394 = 395;
  localparam retro_main_b1_S395 = 396;
  localparam retro_main_b1_S396 = 397;
  localparam retro_main_b1_S397 = 398;
  localparam retro_main_b1_S398 = 399;
  localparam retro_main_b1_S399 = 400;
  localparam retro_main_b1_S400 = 401;
  localparam retro_main_b1_S401 = 402;
  localparam retro_main_b1_S402 = 403;
  localparam retro_main_b1_S403 = 404;
  localparam retro_main_b1_S404 = 405;
  localparam retro_main_b1_S405 = 406;
  localparam retro_main_b1_S406 = 407;
  localparam retro_main_b1_S407 = 408;
  localparam retro_main_b1_S408 = 409;
  localparam retro_main_b1_S409 = 410;
  localparam retro_main_b1_S410 = 411;
  localparam retro_main_b1_S411 = 412;
  localparam retro_main_b1_S412 = 413;
  localparam retro_main_b1_S413 = 414;
  localparam retro_main_b1_S414 = 415;
  localparam retro_main_b1_S415 = 416;
  localparam retro_main_b1_S416 = 417;
  localparam retro_main_b1_S417 = 418;
  localparam retro_main_b1_S418 = 419;
  localparam retro_main_b1_S419 = 420;
  localparam retro_main_b1_S420 = 421;
  localparam retro_main_b1_S421 = 422;
  localparam retro_main_b1_S422 = 423;
  localparam retro_main_b1_S423 = 424;
  localparam retro_main_b1_S424 = 425;
  localparam retro_main_b1_S425 = 426;
  localparam retro_main_b1_S426 = 427;
  localparam retro_main_b1_S427 = 428;
  localparam retro_main_b1_S428 = 429;
  localparam retro_main_b1_S429 = 430;
  localparam retro_main_b1_S430 = 431;
  localparam retro_main_b1_S431 = 432;
  localparam retro_main_b1_S432 = 433;
  localparam retro_main_b1_S433 = 434;
  localparam retro_main_b1_S434 = 435;
  localparam retro_main_b1_S435 = 436;
  localparam retro_main_b1_S436 = 437;
  localparam retro_main_b1_S437 = 438;
  localparam retro_main_b1_S438 = 439;
  localparam retro_main_b1_S439 = 440;
  localparam retro_main_b1_S440 = 441;
  localparam retro_main_b1_S441 = 442;
  localparam retro_main_b1_S442 = 443;
  localparam retro_main_b1_S443 = 444;
  localparam retro_main_b1_S444 = 445;
  localparam retro_main_b1_S445 = 446;
  localparam retro_main_b1_S446 = 447;
  localparam retro_main_b1_S447 = 448;
  localparam retro_main_b1_S448 = 449;
  localparam retro_main_b1_S449 = 450;
  localparam retro_main_b1_S450 = 451;
  localparam retro_main_b1_S451 = 452;
  localparam retro_main_b1_S452 = 453;
  localparam retro_main_b1_S453 = 454;
  localparam retro_main_b1_S454 = 455;
  localparam retro_main_b1_S455 = 456;
  localparam retro_main_b1_S456 = 457;
  localparam retro_main_b1_S457 = 458;
  localparam retro_main_b1_S458 = 459;
  localparam retro_main_b1_S459 = 460;
  localparam retro_main_b1_S460 = 461;
  localparam retro_main_b1_S461 = 462;
  localparam retro_main_b1_S462 = 463;
  localparam retro_main_b1_S463 = 464;
  localparam retro_main_b1_S464 = 465;
  localparam retro_main_b1_S465 = 466;
  localparam retro_main_b1_S466 = 467;
  localparam retro_main_b1_S467 = 468;
  localparam retro_main_b1_S468 = 469;
  localparam retro_main_b1_S469 = 470;
  localparam retro_main_b1_S470 = 471;
  localparam retro_main_b1_S471 = 472;
  localparam retro_main_b1_S472 = 473;
  localparam retro_main_b1_S473 = 474;
  localparam retro_main_b1_S474 = 475;
  localparam retro_main_b1_S475 = 476;
  localparam retro_main_b1_S476 = 477;
  localparam retro_main_b1_S477 = 478;
  localparam retro_main_b1_S478 = 479;
  localparam retro_main_b1_S479 = 480;
  localparam retro_main_b1_S480 = 481;
  localparam retro_main_b1_S481 = 482;
  localparam retro_main_b1_S482 = 483;
  localparam retro_main_b1_S483 = 484;
  localparam retro_main_b1_S484 = 485;
  localparam retro_main_b1_S485 = 486;
  localparam retro_main_b1_S486 = 487;
  localparam retro_main_b1_S487 = 488;
  localparam retro_main_b1_S488 = 489;
  localparam retro_main_b1_S489 = 490;
  localparam retro_main_b1_S490 = 491;
  localparam retro_main_b1_S491 = 492;
  localparam retro_main_b1_S492 = 493;
  localparam retro_main_b1_S493 = 494;
  localparam retro_main_b1_S494 = 495;
  localparam retro_main_b1_S495 = 496;
  localparam retro_main_b1_S496 = 497;
  localparam retro_main_b1_S497 = 498;
  localparam retro_main_b1_S498 = 499;
  localparam retro_main_b1_S499 = 500;
  localparam retro_main_b1_S500 = 501;
  localparam retro_main_b1_S501 = 502;
  localparam retro_main_b1_S502 = 503;
  localparam retro_main_b1_S503 = 504;
  localparam retro_main_b1_S504 = 505;
  localparam retro_main_b1_S505 = 506;
  localparam retro_main_b1_S506 = 507;
  localparam retro_main_b1_S507 = 508;
  localparam retro_main_b1_S508 = 509;
  localparam retro_main_b1_S509 = 510;
  localparam retro_main_b1_S510 = 511;
  localparam retro_main_b1_S511 = 512;
  localparam retro_main_b1_S512 = 513;
  localparam retro_main_b1_S513 = 514;
  localparam retro_main_b1_S514 = 515;
  localparam retro_main_b1_S515 = 516;
  localparam retro_main_b1_S516 = 517;
  localparam retro_main_b1_S517 = 518;
  localparam retro_main_b1_S518 = 519;
  localparam retro_main_b1_S519 = 520;
  localparam retro_main_b1_S520 = 521;
  localparam retro_main_b1_S521 = 522;
  localparam retro_main_b1_S522 = 523;
  localparam retro_main_b1_S523 = 524;
  localparam retro_main_b1_S524 = 525;
  localparam retro_main_b1_S525 = 526;
  localparam retro_main_b1_S526 = 527;
  localparam retro_main_b1_S527 = 528;
  localparam retro_main_b1_S528 = 529;
  localparam retro_main_b1_S529 = 530;
  localparam retro_main_b1_S530 = 531;
  localparam retro_main_b1_S531 = 532;
  localparam retro_main_b1_S532 = 533;
  localparam retro_main_b1_S533 = 534;
  localparam retro_main_b1_S534 = 535;
  localparam retro_main_b1_S535 = 536;
  localparam retro_main_b1_S536 = 537;
  localparam retro_main_b1_S537 = 538;
  localparam retro_main_b1_S538 = 539;
  localparam retro_main_b1_S539 = 540;
  localparam retro_main_b1_S540 = 541;
  localparam retro_main_b1_S541 = 542;
  localparam retro_main_b1_S542 = 543;
  localparam retro_main_b1_S543 = 544;
  localparam retro_main_b1_S544 = 545;
  localparam retro_main_b1_S545 = 546;
  localparam retro_main_b1_S546 = 547;
  localparam retro_main_b1_S547 = 548;
  localparam retro_main_b1_S548 = 549;
  localparam retro_main_b1_S549 = 550;
  localparam retro_main_b1_S550 = 551;
  localparam retro_main_b1_S551 = 552;
  localparam retro_main_b1_S552 = 553;
  localparam retro_main_b1_S553 = 554;
  localparam retro_main_b1_S554 = 555;
  localparam retro_main_b1_S555 = 556;
  localparam retro_main_b1_S556 = 557;
  localparam retro_main_b1_S557 = 558;
  localparam retro_main_b1_S558 = 559;
  localparam retro_main_b1_S559 = 560;
  localparam retro_main_b1_S560 = 561;
  localparam retro_main_b1_S561 = 562;
  localparam retro_main_b1_S562 = 563;
  localparam retro_main_b1_S563 = 564;
  localparam retro_main_b1_S564 = 565;
  localparam retro_main_b1_S565 = 566;
  localparam retro_main_b1_S566 = 567;
  localparam retro_main_b1_S567 = 568;
  localparam retro_main_b1_S568 = 569;
  localparam retro_main_b1_S569 = 570;
  localparam retro_main_b1_S570 = 571;
  localparam retro_main_b1_S571 = 572;
  localparam retro_main_b1_S572 = 573;
  localparam retro_main_b1_S573 = 574;
  localparam retro_main_b1_S574 = 575;
  localparam retro_main_b1_S575 = 576;
  localparam retro_main_b1_S576 = 577;
  localparam retro_main_b1_S577 = 578;
  localparam retro_main_b1_S578 = 579;
  localparam retro_main_b1_S579 = 580;
  localparam retro_main_b1_S580 = 581;
  localparam retro_main_b1_S581 = 582;
  localparam retro_main_b1_S582 = 583;
  localparam retro_main_b1_S583 = 584;
  localparam retro_main_b1_S584 = 585;
  localparam retro_main_b1_S585 = 586;
  localparam retro_main_b1_S586 = 587;
  localparam retro_main_b1_S587 = 588;
  localparam retro_main_b1_S588 = 589;
  localparam retro_main_b1_S589 = 590;
  localparam retro_main_b1_S590 = 591;
  localparam retro_main_b1_S591 = 592;
  localparam retro_main_b1_S592 = 593;
  localparam retro_main_b1_S593 = 594;
  localparam retro_main_b1_S594 = 595;
  localparam retro_main_b1_S595 = 596;
  localparam retro_main_b1_S596 = 597;
  localparam retro_main_b1_S597 = 598;
  localparam retro_main_b1_S598 = 599;
  localparam retro_main_b1_S599 = 600;
  localparam retro_main_b1_S600 = 601;
  localparam retro_main_b1_S601 = 602;
  localparam retro_main_b1_S602 = 603;
  localparam retro_main_b1_S603 = 604;
  localparam retro_main_b1_S604 = 605;
  localparam retro_main_b1_S605 = 606;
  localparam retro_main_b1_S606 = 607;
  localparam retro_main_b1_S607 = 608;
  localparam retro_main_b1_S608 = 609;
  localparam retro_main_b1_S609 = 610;
  localparam retro_main_b1_S610 = 611;
  localparam retro_main_b1_S611 = 612;
  localparam retro_main_b1_S612 = 613;
  localparam retro_main_b1_S613 = 614;
  localparam retro_main_b1_S614 = 615;
  localparam retro_main_b1_S615 = 616;
  localparam retro_main_b1_S616 = 617;
  localparam retro_main_b1_S617 = 618;
  localparam retro_main_b1_S618 = 619;
  localparam retro_main_b1_S619 = 620;
  localparam retro_main_b1_S620 = 621;
  localparam retro_main_b1_S621 = 622;
  localparam retro_main_b1_S622 = 623;
  localparam retro_main_b1_S623 = 624;
  localparam retro_main_b1_S624 = 625;
  localparam retro_main_b1_S625 = 626;
  localparam retro_main_b1_S626 = 627;
  localparam retro_main_b1_S627 = 628;
  localparam retro_main_b1_S628 = 629;
  localparam retro_main_b1_S629 = 630;
  localparam retro_main_b1_S630 = 631;
  localparam retro_main_b1_S631 = 632;
  localparam retro_main_b1_S632 = 633;
  localparam retro_main_b1_S633 = 634;
  localparam retro_main_b1_S634 = 635;
  localparam retro_main_b1_S635 = 636;
  localparam retro_main_b1_S636 = 637;
  localparam retro_main_b1_S637 = 638;
  localparam retro_main_b1_S638 = 639;
  localparam retro_main_b1_S639 = 640;
  localparam retro_main_b1_S640 = 641;
  localparam retro_main_b1_S641 = 642;
  localparam retro_main_b1_S642 = 643;
  localparam retro_main_b1_S643 = 644;
  localparam retro_main_b1_S644 = 645;
  localparam retro_main_b1_S645 = 646;
  localparam retro_main_b1_S646 = 647;
  localparam retro_main_b1_S647 = 648;
  localparam retro_main_b1_S648 = 649;
  localparam retro_main_b1_S649 = 650;
  localparam retro_main_b1_S650 = 651;
  localparam retro_main_b1_S651 = 652;
  localparam retro_main_b1_S652 = 653;
  localparam retro_main_b1_S653 = 654;
  localparam retro_main_b1_S654 = 655;
  localparam retro_main_b1_S655 = 656;
  localparam retro_main_b1_S656 = 657;
  localparam retro_main_b1_S657 = 658;
  localparam retro_main_b1_S658 = 659;
  localparam retro_main_b1_S659 = 660;
  localparam retro_main_b1_S660 = 661;
  localparam retro_main_b1_S661 = 662;
  localparam retro_main_b1_S662 = 663;
  localparam retro_main_b1_S663 = 664;
  localparam retro_main_b1_S664 = 665;
  localparam retro_main_b1_S665 = 666;
  localparam retro_main_b1_S666 = 667;
  localparam retro_main_b1_S667 = 668;
  localparam retro_main_b1_S668 = 669;
  localparam retro_main_b1_S669 = 670;
  localparam retro_main_b1_S670 = 671;
  localparam retro_main_b1_S671 = 672;
  localparam retro_main_b1_S672 = 673;
  localparam retro_main_b1_S673 = 674;
  localparam retro_main_b1_S674 = 675;
  localparam retro_main_b1_S675 = 676;
  localparam retro_main_b1_S676 = 677;
  localparam retro_main_b1_S677 = 678;
  localparam retro_main_b1_S678 = 679;
  localparam retro_main_b1_S679 = 680;
  localparam retro_main_b1_S680 = 681;
  localparam retro_main_b1_S681 = 682;
  localparam retro_main_b1_S682 = 683;
  localparam retro_main_b1_S683 = 684;
  localparam retro_main_b1_S684 = 685;
  localparam retro_main_b1_S685 = 686;
  localparam retro_main_b1_S686 = 687;
  localparam retro_main_b1_S687 = 688;
  localparam retro_main_b1_S688 = 689;
  localparam retro_main_b1_S689 = 690;
  localparam retro_main_b1_S690 = 691;
  localparam retro_main_b1_S691 = 692;
  localparam retro_main_b1_S692 = 693;
  localparam retro_main_b1_S693 = 694;
  localparam retro_main_b1_S694 = 695;
  localparam retro_main_b1_S695 = 696;
  localparam retro_main_b1_S696 = 697;
  localparam retro_main_b1_S697 = 698;
  localparam retro_main_b1_S698 = 699;
  localparam retro_main_b1_S699 = 700;
  localparam retro_main_b1_S700 = 701;
  localparam retro_main_b1_S701 = 702;
  localparam retro_main_b1_S702 = 703;
  localparam retro_main_b1_S703 = 704;
  localparam retro_main_b1_S704 = 705;
  localparam retro_main_b1_S705 = 706;
  localparam retro_main_b1_S706 = 707;
  localparam retro_main_b1_S707 = 708;
  localparam retro_main_b1_S708 = 709;
  localparam retro_main_b1_S709 = 710;
  localparam retro_main_b1_S710 = 711;
  localparam retro_main_b1_S711 = 712;
  localparam retro_main_b1_S712 = 713;
  localparam retro_main_b1_S713 = 714;
  localparam retro_main_b1_S714 = 715;
  localparam retro_main_b1_S715 = 716;
  localparam retro_main_b1_S716 = 717;
  localparam retro_main_b1_S717 = 718;
  localparam retro_main_b1_S718 = 719;
  localparam retro_main_b1_S719 = 720;
  localparam retro_main_b1_S720 = 721;
  localparam retro_main_b1_S721 = 722;
  localparam retro_main_b1_S722 = 723;
  localparam retro_main_b1_S723 = 724;
  localparam retro_main_b1_S724 = 725;
  localparam retro_main_b1_S725 = 726;
  localparam retro_main_b1_S726 = 727;
  localparam retro_main_b1_S727 = 728;
  localparam retro_main_b1_S728 = 729;
  localparam retro_main_b1_S729 = 730;
  localparam retro_main_b1_S730 = 731;
  localparam retro_main_b1_S731 = 732;
  localparam retro_main_b1_S732 = 733;
  localparam retro_main_b1_S733 = 734;
  localparam retro_main_b1_S734 = 735;
  localparam retro_main_b1_S735 = 736;
  localparam retro_main_b1_S736 = 737;
  localparam retro_main_b1_S737 = 738;
  localparam retro_main_b1_S738 = 739;
  localparam retro_main_b1_S739 = 740;
  localparam retro_main_b1_S740 = 741;
  localparam retro_main_b1_S741 = 742;
  localparam retro_main_b1_S742 = 743;
  localparam retro_main_b1_S743 = 744;
  localparam retro_main_b1_S744 = 745;
  localparam retro_main_b1_S745 = 746;
  localparam retro_main_b1_S746 = 747;
  localparam retro_main_b1_S747 = 748;
  localparam retro_main_b1_S748 = 749;
  localparam retro_main_b1_S749 = 750;
  localparam retro_main_b1_S750 = 751;
  localparam retro_main_b1_S751 = 752;
  localparam retro_main_b1_S752 = 753;
  localparam retro_main_b1_S753 = 754;
  localparam retro_main_b1_S754 = 755;
  localparam retro_main_b1_S755 = 756;
  localparam retro_main_b1_S756 = 757;
  localparam retro_main_b1_S757 = 758;
  localparam retro_main_b1_S758 = 759;
  localparam retro_main_b1_S759 = 760;
  localparam retro_main_b1_S760 = 761;
  localparam retro_main_b1_S761 = 762;
  localparam retro_main_b1_S762 = 763;
  localparam retro_main_b1_S763 = 764;
  localparam retro_main_b1_S764 = 765;
  localparam retro_main_b1_S765 = 766;
  localparam retro_main_b1_S766 = 767;
  localparam retro_main_b1_S767 = 768;
  localparam retro_main_b1_S768 = 769;
  localparam retro_main_b1_S769 = 770;
  localparam retro_main_b1_S770 = 771;
  localparam retro_main_b1_S771 = 772;
  localparam retro_main_b1_S772 = 773;
  localparam retro_main_b1_S773 = 774;
  localparam retro_main_b1_S774 = 775;
  localparam retro_main_b1_S775 = 776;
  localparam retro_main_b1_S776 = 777;
  localparam retro_main_b1_S777 = 778;
  localparam retro_main_b1_S778 = 779;
  localparam retro_main_b1_S779 = 780;
  localparam retro_main_b1_S780 = 781;
  localparam retro_main_b1_S781 = 782;
  localparam retro_main_b1_S782 = 783;
  localparam retro_main_b1_S783 = 784;
  localparam retro_main_b1_S784 = 785;
  localparam retro_main_b1_S785 = 786;
  localparam retro_main_b1_S786 = 787;
  localparam retro_main_b1_S787 = 788;
  localparam retro_main_b1_S788 = 789;
  localparam retro_main_b1_S789 = 790;
  localparam retro_main_b1_S790 = 791;
  localparam retro_main_b1_S791 = 792;
  localparam retro_main_b1_S792 = 793;
  localparam retro_main_b1_S793 = 794;
  localparam retro_main_b1_S794 = 795;
  localparam retro_main_b1_S795 = 796;
  localparam retro_main_b1_S796 = 797;
  localparam retro_main_b1_S797 = 798;
  localparam retro_main_b1_S798 = 799;
  localparam retro_main_b1_S799 = 800;
  localparam retro_main_b1_S800 = 801;
  localparam retro_main_b1_S801 = 802;
  localparam retro_main_b1_S802 = 803;
  localparam retro_main_b1_S803 = 804;
  localparam retro_main_b1_S804 = 805;
  localparam retro_main_b1_S805 = 806;
  localparam retro_main_b1_S806 = 807;
  localparam retro_main_b1_S807 = 808;
  localparam retro_main_b1_S808 = 809;
  localparam retro_main_b1_S809 = 810;
  localparam retro_main_b1_S810 = 811;
  localparam retro_main_b1_S811 = 812;
  localparam retro_main_b1_S812 = 813;
  localparam retro_main_b1_S813 = 814;
  localparam retro_main_b1_S814 = 815;
  localparam retro_main_b1_S815 = 816;
  localparam retro_main_b1_S816 = 817;
  localparam retro_main_b1_S817 = 818;
  localparam retro_main_b1_S818 = 819;
  localparam retro_main_b1_S819 = 820;
  localparam retro_main_b1_S820 = 821;
  localparam retro_main_b1_S821 = 822;
  localparam retro_main_b1_S822 = 823;
  localparam retro_main_b1_S823 = 824;
  localparam retro_main_b1_S824 = 825;
  localparam retro_main_b1_S825 = 826;
  localparam retro_main_b1_S826 = 827;
  localparam retro_main_b1_S827 = 828;
  localparam retro_main_b1_S828 = 829;
  localparam retro_main_b1_S829 = 830;
  localparam retro_main_b1_S830 = 831;
  localparam retro_main_b1_S831 = 832;
  localparam retro_main_b1_S832 = 833;
  localparam retro_main_b1_S833 = 834;
  localparam retro_main_b1_S834 = 835;
  localparam retro_main_b1_S835 = 836;
  localparam retro_main_b1_S836 = 837;
  localparam retro_main_b1_S837 = 838;
  localparam retro_main_b1_S838 = 839;
  localparam retro_main_b1_S839 = 840;
  localparam retro_main_b1_S840 = 841;
  localparam retro_main_b1_S841 = 842;
  localparam retro_main_b1_S842 = 843;
  localparam retro_main_b1_S843 = 844;
  localparam retro_main_b1_S844 = 845;
  localparam retro_main_b1_S845 = 846;
  localparam retro_main_b1_S846 = 847;
  localparam retro_main_b1_S847 = 848;
  localparam retro_main_b1_S848 = 849;
  localparam retro_main_b1_S849 = 850;
  localparam retro_main_b1_S850 = 851;
  localparam retro_main_b1_S851 = 852;
  localparam retro_main_b1_S852 = 853;
  localparam retro_main_b1_S853 = 854;
  localparam retro_main_b1_S854 = 855;
  localparam retro_main_b1_S855 = 856;
  localparam retro_main_b1_S856 = 857;
  localparam retro_main_b1_S857 = 858;
  localparam retro_main_b1_S858 = 859;
  localparam retro_main_b1_S859 = 860;
  localparam retro_main_b1_S860 = 861;
  localparam retro_main_b1_S861 = 862;
  localparam retro_main_b1_S862 = 863;
  localparam retro_main_b1_S863 = 864;
  localparam retro_main_b1_S864 = 865;
  localparam retro_main_b1_S865 = 866;
  localparam retro_main_b1_S866 = 867;
  localparam retro_main_b1_S867 = 868;
  localparam retro_main_b1_S868 = 869;
  localparam retro_main_b1_S869 = 870;
  localparam retro_main_b1_S870 = 871;
  localparam retro_main_b1_S871 = 872;
  localparam retro_main_b1_S872 = 873;
  localparam retro_main_b1_S873 = 874;
  localparam retro_main_b1_S874 = 875;
  localparam retro_main_b1_S875 = 876;
  localparam retro_main_b1_S876 = 877;
  localparam retro_main_b1_S877 = 878;
  localparam retro_main_b1_S878 = 879;
  localparam retro_main_b1_S879 = 880;
  localparam retro_main_b1_S880 = 881;
  localparam retro_main_b1_S881 = 882;
  localparam retro_main_b1_S882 = 883;
  localparam retro_main_b1_S883 = 884;
  localparam retro_main_b1_S884 = 885;
  localparam retro_main_b1_S885 = 886;
  localparam retro_main_b1_S886 = 887;
  localparam retro_main_b1_S887 = 888;
  localparam retro_main_b1_S888 = 889;
  localparam retro_main_b1_S889 = 890;
  localparam retro_main_b1_S890 = 891;
  localparam retro_main_b1_S891 = 892;
  localparam retro_main_b1_S892 = 893;
  localparam retro_main_b1_S893 = 894;
  localparam retro_main_b1_S894 = 895;
  localparam retro_main_b1_S895 = 896;
  localparam retro_main_b1_S896 = 897;
  localparam retro_main_b1_S897 = 898;
  localparam retro_main_b1_S898 = 899;
  localparam retro_main_b1_S899 = 900;
  localparam retro_main_b1_S900 = 901;
  localparam retro_main_b1_S901 = 902;
  localparam retro_main_b1_S902 = 903;
  localparam retro_main_b1_S903 = 904;
  localparam retro_main_b1_S904 = 905;
  localparam retro_main_b1_S905 = 906;
  localparam retro_main_b1_S906 = 907;
  localparam retro_main_b1_S907 = 908;
  localparam retro_main_b1_S908 = 909;
  localparam retro_main_b1_S909 = 910;
  localparam retro_main_b1_S910 = 911;
  localparam retro_main_b1_S911 = 912;
  localparam retro_main_b1_S912 = 913;
  localparam retro_main_b1_S913 = 914;
  localparam retro_main_b1_S914 = 915;
  localparam retro_main_b1_S915 = 916;
  localparam retro_main_b1_S916 = 917;
  localparam retro_main_b1_S917 = 918;
  localparam retro_main_b1_S918 = 919;
  localparam retro_main_b1_S919 = 920;
  localparam retro_main_b1_S920 = 921;
  localparam retro_main_b1_S921 = 922;
  localparam retro_main_b1_S922 = 923;
  localparam retro_main_b1_S923 = 924;
  localparam retro_main_b1_S924 = 925;
  localparam retro_main_b1_S925 = 926;
  localparam retro_main_b1_S926 = 927;
  localparam retro_main_b1_S927 = 928;
  localparam retro_main_b1_S928 = 929;
  localparam retro_main_b1_S929 = 930;
  localparam retro_main_b1_S930 = 931;
  localparam retro_main_b1_S931 = 932;
  localparam retro_main_b1_S932 = 933;
  localparam retro_main_b1_S933 = 934;
  localparam retro_main_b1_S934 = 935;
  localparam retro_main_b1_S935 = 936;
  localparam retro_main_b1_S936 = 937;
  localparam retro_main_b1_S937 = 938;
  localparam retro_main_b1_S938 = 939;
  localparam retro_main_b1_S939 = 940;
  localparam retro_main_b1_S940 = 941;
  localparam retro_main_b1_S941 = 942;
  localparam retro_main_b1_S942 = 943;
  localparam retro_main_b1_S943 = 944;
  localparam retro_main_b1_S944 = 945;
  localparam retro_main_b1_S945 = 946;
  localparam retro_main_b1_S946 = 947;
  localparam retro_main_b1_S947 = 948;
  localparam retro_main_b1_S948 = 949;
  localparam retro_main_b1_S949 = 950;
  localparam retro_main_b1_S950 = 951;
  localparam retro_main_b1_S951 = 952;
  localparam retro_main_b1_S952 = 953;
  localparam retro_main_b1_S953 = 954;
  localparam retro_main_b1_S954 = 955;
  localparam retro_main_b1_S955 = 956;
  localparam retro_main_b1_S956 = 957;
  localparam retro_main_b1_S957 = 958;
  localparam retro_main_b1_S958 = 959;
  localparam retro_main_b1_S959 = 960;
  localparam retro_main_b1_S960 = 961;
  localparam retro_main_b1_S961 = 962;
  localparam retro_main_b1_S962 = 963;
  localparam retro_main_b1_S963 = 964;
  localparam retro_main_b1_S964 = 965;
  localparam retro_main_b1_S965 = 966;
  localparam retro_main_b1_S966 = 967;
  localparam retro_main_b1_S967 = 968;
  localparam retro_main_b1_S968 = 969;
  localparam retro_main_b1_S969 = 970;
  localparam retro_main_b1_S970 = 971;
  localparam retro_main_b1_S971 = 972;
  localparam retro_main_b1_S972 = 973;
  localparam retro_main_b1_S973 = 974;
  localparam retro_main_b1_S974 = 975;
  localparam retro_main_b1_S975 = 976;
  localparam retro_main_b1_S976 = 977;
  localparam retro_main_b1_S977 = 978;
  localparam retro_main_b1_S978 = 979;
  localparam retro_main_b1_S979 = 980;
  localparam retro_main_b1_S980 = 981;
  localparam retro_main_b1_S981 = 982;
  localparam retro_main_b1_S982 = 983;
  localparam retro_main_b1_S983 = 984;
  localparam retro_main_b1_S984 = 985;
  localparam retro_main_b1_S985 = 986;
  localparam retro_main_b1_S986 = 987;
  localparam retro_main_b1_S987 = 988;
  localparam retro_main_b1_S988 = 989;
  localparam retro_main_b1_S989 = 990;
  localparam retro_main_b1_S990 = 991;
  localparam retro_main_b1_S991 = 992;
  localparam retro_main_b1_S992 = 993;
  localparam retro_main_b1_S993 = 994;
  localparam retro_main_b1_S994 = 995;
  localparam retro_main_b1_S995 = 996;
  localparam retro_main_b1_S996 = 997;
  localparam retro_main_b1_S997 = 998;
  localparam retro_main_b1_S998 = 999;
  localparam retro_main_b1_S999 = 1000;
  localparam retro_main_b1_S1000 = 1001;
  localparam retro_main_b1_S1001 = 1002;
  localparam retro_main_b1_S1002 = 1003;
  localparam retro_main_b1_S1003 = 1004;
  localparam retro_main_b1_S1004 = 1005;
  localparam retro_main_b1_S1005 = 1006;
  localparam retro_main_b1_S1006 = 1007;
  localparam retro_main_b1_S1007 = 1008;
  localparam retro_main_b1_S1008 = 1009;
  localparam retro_main_b1_S1009 = 1010;
  localparam retro_main_b1_S1010 = 1011;
  localparam retro_main_b1_S1011 = 1012;
  localparam retro_main_b1_S1012 = 1013;
  localparam retro_main_b1_S1013 = 1014;
  localparam retro_main_b1_S1014 = 1015;
  localparam retro_main_b1_S1015 = 1016;
  localparam retro_main_b1_S1016 = 1017;
  localparam retro_main_b1_S1017 = 1018;
  localparam retro_main_b1_S1018 = 1019;
  localparam retro_main_b1_S1019 = 1020;
  localparam retro_main_b1_S1020 = 1021;
  localparam retro_main_b1_S1021 = 1022;
  localparam retro_main_b1_S1022 = 1023;
  localparam retro_main_b1_S1023 = 1024;
  localparam retro_main_b1_S1024 = 1025;
  localparam retro_main_whileelse200_FINISH = 1026;
  localparam retro_main_L1_while2_S0 = 1027;
  localparam retro_main_L1_whilebody3_S0 = 1028;
  localparam retro_main_L1_whilebody3_S1 = 1029;
  localparam retro_main_L1_whilebody3_S2 = 1030;
  localparam retro_main_L1_whilebody3_S3 = 1031;
  localparam retro_main_L1_whilebody3_S4 = 1032;
  localparam retro_main_L1_ifthen4_S0 = 1033;
  localparam retro_main_L1_ifelse197_S0 = 1034;
  localparam retro_main_L1_ifelse197_S1 = 1035;
  localparam retro_main_L1_ifelse197_S2 = 1036;
  localparam retro_main_L1_ifelse197_S3 = 1037;
  localparam retro_main_L1_ifthen11_S0 = 1038;
  localparam retro_main_L1_ifthen11_S1 = 1039;
  localparam retro_main_L1_ifthen11_S2 = 1040;
  localparam retro_main_L1_ifthen11_S3 = 1041;
  localparam retro_main_L1_ifthen15_S0 = 1042;
  localparam retro_main_L1_ifthen15_S1 = 1043;
  localparam retro_main_L1_ifthen19_S0 = 1044;
  localparam retro_main_L1_ifthen19_S1 = 1045;
  localparam retro_main_L1_ifthen19_S2 = 1046;
  localparam retro_main_L1_ifthen19_S3 = 1047;
  localparam retro_main_L1_ifthen23_S0 = 1048;
  localparam retro_main_L1_ifthen27_S0 = 1049;
  localparam retro_main_L1_ifthen27_S1 = 1050;
  localparam retro_main_L1_ifthen27_S2 = 1051;
  localparam retro_main_L1_ifthen27_S3 = 1052;
  localparam retro_main_L1_ifthen31_S0 = 1053;
  localparam retro_main_L1_ifthen31_S1 = 1054;
  localparam retro_main_L1_ifthen31_S2 = 1055;
  localparam retro_main_L1_ifthen31_S3 = 1056;
  localparam retro_main_L1_ifthen35_S0 = 1057;
  localparam retro_main_L1_ifthen44_S0 = 1058;
  localparam retro_main_L1_ifthen44_S1 = 1059;
  localparam retro_main_L1_ifthen44_S2 = 1060;
  localparam retro_main_L1_ifthen44_S3 = 1061;
  localparam retro_main_L1_ifthen48_S0 = 1062;
  localparam retro_main_L1_ifthen48_S1 = 1063;
  localparam retro_main_L1_ifthen48_S2 = 1064;
  localparam retro_main_L1_ifthen48_S3 = 1065;
  localparam retro_main_L1_ifthen52_S0 = 1066;
  localparam retro_main_L1_ifthen52_S1 = 1067;
  localparam retro_main_L1_ifthen52_S2 = 1068;
  localparam retro_main_L1_ifthen52_S3 = 1069;
  localparam retro_main_L1_ifthen52_S4 = 1070;
  localparam retro_main_L1_ifthen61_S0 = 1071;
  localparam retro_main_L1_ifthen61_S1 = 1072;
  localparam retro_main_L1_ifthen61_S2 = 1073;
  localparam retro_main_L1_ifthen61_S3 = 1074;
  localparam retro_main_L1_ifthen61_S4 = 1075;
  localparam retro_main_L1_ifthen70_S0 = 1076;
  localparam retro_main_L1_ifthen70_S1 = 1077;
  localparam retro_main_L1_ifthen70_S2 = 1078;
  localparam retro_main_L1_ifthen70_S3 = 1079;
  localparam retro_main_L1_ifthen70_S4 = 1080;
  localparam retro_main_L1_ifthen79_S0 = 1081;
  localparam retro_main_L1_ifthen79_S1 = 1082;
  localparam retro_main_L1_ifthen79_S2 = 1083;
  localparam retro_main_L1_ifthen79_S3 = 1084;
  localparam retro_main_L1_ifthen79_S4 = 1085;
  localparam retro_main_L1_ifthen88_S0 = 1086;
  localparam retro_main_L1_ifthen88_S1 = 1087;
  localparam retro_main_L1_ifthen88_S2 = 1088;
  localparam retro_main_L1_ifthen88_S3 = 1089;
  localparam retro_main_L1_ifthen92_S0 = 1090;
  localparam retro_main_L1_ifthen92_S1 = 1091;
  localparam retro_main_L1_ifthen92_S2 = 1092;
  localparam retro_main_L1_ifthen92_S3 = 1093;
  localparam retro_main_L1_ifthen92_S4 = 1094;
  localparam retro_main_L1_ifthen96_S0 = 1095;
  localparam retro_main_L1_ifthen96_S1 = 1096;
  localparam retro_main_L1_ifthen96_S2 = 1097;
  localparam retro_main_L1_ifthen96_S3 = 1098;
  localparam retro_main_L1_ifthen100_S0 = 1099;
  localparam retro_main_L1_ifthen100_S1 = 1100;
  localparam retro_main_L1_ifthen100_S2 = 1101;
  localparam retro_main_L1_ifthen100_S3 = 1102;
  localparam retro_main_L1_ifthen104_S0 = 1103;
  localparam retro_main_L1_ifthen104_S1 = 1104;
  localparam retro_main_L1_ifthen104_S2 = 1105;
  localparam retro_main_L1_ifthen104_S3 = 1106;
  localparam retro_main_L1_ifthen108_S0 = 1107;
  localparam retro_main_L1_ifthen108_S1 = 1108;
  localparam retro_main_L1_ifthen112_S0 = 1109;
  localparam retro_main_L1_ifthen112_S1 = 1110;
  localparam retro_main_L1_ifthen112_S2 = 1111;
  localparam retro_main_L1_ifthen112_S3 = 1112;
  localparam retro_main_L1_ifthen116_S0 = 1113;
  localparam retro_main_L1_ifthen116_S1 = 1114;
  localparam retro_main_L1_ifthen116_S2 = 1115;
  localparam retro_main_L1_ifthen116_S3 = 1116;
  localparam retro_main_L1_ifthen120_S0 = 1117;
  localparam retro_main_L1_ifthen120_S1 = 1118;
  localparam retro_main_L1_ifthen120_S2 = 1119;
  localparam retro_main_L1_ifthen120_S3 = 1120;
  localparam retro_main_L1_ifthen124_S0 = 1121;
  localparam retro_main_L1_ifthen124_S1 = 1122;
  localparam retro_main_L1_ifthen124_S2 = 1123;
  localparam retro_main_L1_ifthen124_S3 = 1124;
  localparam retro_main_L1_ifthen128_S0 = 1125;
  localparam retro_main_L1_ifthen128_S1 = 1126;
  localparam retro_main_L1_ifthen128_S2 = 1127;
  localparam retro_main_L1_ifthen128_S3 = 1128;
  localparam retro_main_L1_ifthen132_S0 = 1129;
  localparam retro_main_L1_ifthen141_S0 = 1130;
  localparam retro_main_L1_ifthen145_S0 = 1131;
  localparam retro_main_L1_ifthen149_S0 = 1132;
  localparam retro_main_L1_ifthen149_S1 = 1133;
  localparam retro_main_L1_ifthen153_S0 = 1134;
  localparam retro_main_L1_ifthen153_S1 = 1135;
  localparam retro_main_L1_ifthen153_S2 = 1136;
  localparam retro_main_L1_ifthen153_S3 = 1137;
  localparam retro_main_L1_ifthen153_S4 = 1138;
  localparam retro_main_L1_ifthen157_S0 = 1139;
  localparam retro_main_L1_ifthen157_S1 = 1140;
  localparam retro_main_L1_ifthen38_S0 = 1141;
  localparam retro_main_L1_ifthen38_S1 = 1142;
  localparam retro_main_L1_ifthen38_S2 = 1143;
  localparam retro_main_L1_ifthen38_S3 = 1144;
  localparam retro_main_L1_ifelse41_S0 = 1145;
  localparam retro_main_L1_ifelse41_S1 = 1146;
  localparam retro_main_L1_ifelse41_S2 = 1147;
  localparam retro_main_L1_ifelse41_S3 = 1148;
  localparam retro_main_L1_ifthen55_S0 = 1149;
  localparam retro_main_L1_ifthen55_S1 = 1150;
  localparam retro_main_L1_ifthen55_S2 = 1151;
  localparam retro_main_L1_ifthen55_S3 = 1152;
  localparam retro_main_L1_ifthen64_S0 = 1153;
  localparam retro_main_L1_ifthen64_S1 = 1154;
  localparam retro_main_L1_ifthen64_S2 = 1155;
  localparam retro_main_L1_ifthen64_S3 = 1156;
  localparam retro_main_L1_ifthen73_S0 = 1157;
  localparam retro_main_L1_ifthen73_S1 = 1158;
  localparam retro_main_L1_ifthen73_S2 = 1159;
  localparam retro_main_L1_ifthen73_S3 = 1160;
  localparam retro_main_L1_ifthen82_S0 = 1161;
  localparam retro_main_L1_ifthen82_S1 = 1162;
  localparam retro_main_L1_ifthen82_S2 = 1163;
  localparam retro_main_L1_ifthen82_S3 = 1164;
  localparam retro_main_L1_ifthen135_S0 = 1165;
  localparam retro_main_L1_ifthen135_S1 = 1166;
  localparam retro_main_L1_ifthen135_S2 = 1167;
  localparam retro_main_L1_ifthen135_S3 = 1168;
  localparam retro_main_L1_ifthen160_S0 = 1169;
  localparam retro_main_L1_ifthen160_S1 = 1170;
  localparam retro_main_L1_b603_S0 = 1171;
  localparam retro_main_L1_b604_S0 = 1172;
  localparam retro_main_L1_b605_S0 = 1173;
  localparam retro_main_L1_b606_S0 = 1174;
  localparam retro_main_L1_ifthen424_S0 = 1175;
  localparam retro_main_L1_ifthen395_S0 = 1176;
  localparam retro_main_L1_exit396_S0 = 1177;
  localparam retro_main_L1_exit396_S1 = 1178;
  localparam retro_main_L1_whileexit429_S0 = 1179;
  localparam retro_main_L1_whileexit429_S1 = 1180;
  localparam retro_main_L1_whileexit434_S0 = 1181;
  localparam retro_main_L1_whileexit434_S1 = 1182;
  localparam retro_main_L1_whileexit434_S2 = 1183;
  localparam retro_main_L1_whileexit434_S3 = 1184;
  localparam retro_main_L1_ifthen401_S0 = 1185;
  localparam retro_main_L1_exit402_S0 = 1186;
  localparam retro_main_L1_exit402_S1 = 1187;
  localparam retro_main_L1_whileexit439_S0 = 1188;
  localparam retro_main_L1_whileexit439_S1 = 1189;
  localparam retro_main_L1_whileexit439_S2 = 1190;
  localparam retro_main_L1_ifthen442_S0 = 1191;
  localparam retro_main_L1_ifthen442_S1 = 1192;
  localparam retro_main_L1_forelse409_S0 = 1193;
  localparam retro_main_L1_forelse409_S2 = 1194;
  localparam retro_main_L1_b443_S0 = 1195;
  localparam retro_main_L1_b443_S1 = 1196;
  localparam retro_main_L1_ifthen444_S0 = 1197;
  localparam retro_main_L1_ifthen445_S0 = 1198;
  localparam retro_main_L1_ifelse594_S0 = 1199;
  localparam retro_main_L1_ifelse594_S1 = 1200;
  localparam retro_main_L1_ifelse594_S2 = 1201;
  localparam retro_main_L1_ifelse594_S3 = 1202;
  localparam retro_main_L1_ifthen446_S0 = 1203;
  localparam retro_main_L1_ifthen446_S1 = 1204;
  localparam retro_main_L1_ifthen446_S2 = 1205;
  localparam retro_main_L1_ifthen446_S3 = 1206;
  localparam retro_main_L1_ifelse569_S0 = 1207;
  localparam retro_main_L1_ifelse569_S1 = 1208;
  localparam retro_main_L1_ifelse569_S2 = 1209;
  localparam retro_main_L1_ifelse569_S3 = 1210;
  localparam retro_main_L1_whileexit455_S0 = 1211;
  localparam retro_main_L1_whileexit455_S1 = 1212;
  localparam retro_main_L1_whileexit455_S2 = 1213;
  localparam retro_main_L1_whileexit578_S0 = 1214;
  localparam retro_main_L1_whileexit578_S1 = 1215;
  localparam retro_main_L1_whileexit578_S2 = 1216;
  localparam retro_main_L1_whileexit460_S0 = 1217;
  localparam retro_main_L1_whileexit460_S1 = 1218;
  localparam retro_main_L1_whileexit583_S0 = 1219;
  localparam retro_main_L1_whileexit583_S1 = 1220;
  localparam retro_main_L1_whileexit472_S0 = 1221;
  localparam retro_main_L1_whileexit472_S1 = 1222;
  localparam retro_main_L1_whileexit472_S2 = 1223;
  localparam retro_main_L1_whileexit477_S0 = 1224;
  localparam retro_main_L1_whileexit477_S1 = 1225;
  localparam retro_main_L1_whileexit489_S0 = 1226;
  localparam retro_main_L1_whileexit489_S1 = 1227;
  localparam retro_main_L1_whileexit489_S2 = 1228;
  localparam retro_main_L1_whileexit494_S0 = 1229;
  localparam retro_main_L1_whileexit494_S1 = 1230;
  localparam retro_main_L1_b502_S0 = 1231;
  localparam retro_main_L1_whileexit507_S0 = 1232;
  localparam retro_main_L1_whileexit507_S1 = 1233;
  localparam retro_main_L1_whileexit512_S0 = 1234;
  localparam retro_main_L1_whileexit512_S1 = 1235;
  localparam retro_main_L1_whileexit517_S0 = 1236;
  localparam retro_main_L1_whileexit517_S1 = 1237;
  localparam retro_main_L1_b520_S0 = 1238;
  localparam retro_main_L1_b520_S1 = 1239;
  localparam retro_main_L1_ifthen521_S0 = 1240;
  localparam retro_main_L1_ifthen521_S1 = 1241;
  localparam retro_main_L1_b522_S0 = 1242;
  localparam retro_main_L1_b522_S1 = 1243;
  localparam retro_main_L1_ifthen523_S0 = 1244;
  localparam retro_main_L1_ifthen523_S1 = 1245;
  localparam retro_main_L1_b524_S0 = 1246;
  localparam retro_main_L1_b524_S1 = 1247;
  localparam retro_main_L1_ifthen525_S0 = 1248;
  localparam retro_main_L1_ifthen525_S1 = 1249;
  localparam retro_main_L1_ifthen551_S0 = 1250;
  localparam retro_main_L1_ifthen551_S1 = 1251;
  localparam retro_main_L1_ifthen552_S0 = 1252;
  localparam retro_main_L1_ifthen552_S1 = 1253;
  localparam retro_main_L1_ifthen553_S0 = 1254;
  localparam retro_main_L1_ifthen553_S1 = 1255;
  localparam retro_main_L1_ifthen554_S0 = 1256;
  localparam retro_main_L1_ifthen554_S1 = 1257;
  localparam retro_main_L1_ifthen555_S0 = 1258;
  localparam retro_main_L1_ifthen555_S1 = 1259;
  localparam retro_main_L1_ifthen556_S0 = 1260;
  localparam retro_main_L1_ifthen556_S1 = 1261;
  localparam retro_main_L1_b526_S0 = 1262;
  localparam retro_main_L1_b526_S1 = 1263;
  localparam retro_main_L1_ifthen527_S0 = 1264;
  localparam retro_main_L1_ifthen527_S1 = 1265;
  localparam retro_main_L1_b528_S0 = 1266;
  localparam retro_main_L1_b528_S1 = 1267;
  localparam retro_main_L1_ifthen529_S0 = 1268;
  localparam retro_main_L1_ifthen529_S1 = 1269;
  localparam retro_main_L1_ifthen533_S0 = 1270;
  localparam retro_main_L1_ifthen533_S1 = 1271;
  localparam retro_main_L1_ifthen534_S0 = 1272;
  localparam retro_main_L1_ifthen534_S1 = 1273;
  localparam retro_main_L1_ifthen535_S0 = 1274;
  localparam retro_main_L1_ifthen535_S1 = 1275;
  localparam retro_main_L1_ifthen536_S0 = 1276;
  localparam retro_main_L1_ifthen536_S1 = 1277;
  localparam retro_main_L1_ifthen539_S0 = 1278;
  localparam retro_main_L1_ifthen539_S1 = 1279;
  localparam retro_main_L1_ifthen542_S0 = 1280;
  localparam retro_main_L1_ifthen542_S1 = 1281;
  localparam retro_main_L1_ifthen543_S0 = 1282;
  localparam retro_main_L1_ifthen543_S1 = 1283;
  localparam retro_main_L1_ifthen544_S0 = 1284;
  localparam retro_main_L1_ifthen544_S1 = 1285;
  localparam retro_main_L1_ifthen545_S0 = 1286;
  localparam retro_main_L1_ifthen545_S1 = 1287;
  localparam retro_main_L1_ifthen546_S0 = 1288;
  localparam retro_main_L1_ifthen546_S1 = 1289;
  localparam retro_main_L1_ifthen547_S0 = 1290;
  localparam retro_main_L1_ifthen547_S1 = 1291;
  localparam retro_main_L1_ifthen548_S0 = 1292;
  localparam retro_main_L1_ifthen548_S1 = 1293;
  localparam retro_main_L1_ifthen549_S0 = 1294;
  localparam retro_main_L1_ifthen549_S1 = 1295;
  localparam retro_main_L1_ifthen550_S0 = 1296;
  localparam retro_main_L1_ifthen550_S1 = 1297;
  localparam retro_main_L1_b530_S0 = 1298;
  localparam retro_main_L1_b530_S1 = 1299;
  localparam retro_main_L1_ifthen531_S0 = 1300;
  localparam retro_main_L1_ifthen531_S1 = 1301;
  localparam retro_main_L1_b532_S0 = 1302;
  localparam retro_main_L1_b198_S0 = 1303;
  localparam retro_main_L1_b198_S1 = 1304;
  localparam retro_main_L2_while427_S0 = 1305;
  localparam retro_main_L2_while427_S1 = 1306;
  localparam retro_main_L2_while427_S2 = 1307;
  localparam retro_main_L2_while427_S3 = 1308;
  localparam retro_main_L2_ifelse601_S0 = 1309;
  localparam retro_main_L3_while432_S0 = 1310;
  localparam retro_main_L3_while432_S1 = 1311;
  localparam retro_main_L3_while432_S2 = 1312;
  localparam retro_main_L3_while432_S3 = 1313;
  localparam retro_main_L3_ifelse600_S0 = 1314;
  localparam retro_main_L4_while437_S0 = 1315;
  localparam retro_main_L4_while437_S1 = 1316;
  localparam retro_main_L4_while437_S2 = 1317;
  localparam retro_main_L4_while437_S3 = 1318;
  localparam retro_main_L4_ifelse599_S0 = 1319;
  localparam retro_main_L5_while576_S0 = 1320;
  localparam retro_main_L5_while576_S1 = 1321;
  localparam retro_main_L5_while576_S2 = 1322;
  localparam retro_main_L5_while576_S3 = 1323;
  localparam retro_main_L5_ifelse593_S0 = 1324;
  localparam retro_main_L6_while581_S0 = 1325;
  localparam retro_main_L6_while581_S1 = 1326;
  localparam retro_main_L6_while581_S2 = 1327;
  localparam retro_main_L6_while581_S3 = 1328;
  localparam retro_main_L6_ifelse592_S0 = 1329;
  localparam retro_main_L7_while586_S0 = 1330;
  localparam retro_main_L7_while586_S1 = 1331;
  localparam retro_main_L7_while586_S2 = 1332;
  localparam retro_main_L7_while586_S3 = 1333;
  localparam retro_main_L7_ifelse591_S0 = 1334;
  localparam retro_main_L8_while453_S0 = 1335;
  localparam retro_main_L8_while453_S1 = 1336;
  localparam retro_main_L8_while453_S2 = 1337;
  localparam retro_main_L8_while453_S3 = 1338;
  localparam retro_main_L8_ifelse568_S0 = 1339;
  localparam retro_main_L9_while458_S0 = 1340;
  localparam retro_main_L9_while458_S1 = 1341;
  localparam retro_main_L9_while458_S2 = 1342;
  localparam retro_main_L9_while458_S3 = 1343;
  localparam retro_main_L9_ifelse567_S0 = 1344;
  localparam retro_main_L10_while463_S0 = 1345;
  localparam retro_main_L10_while463_S1 = 1346;
  localparam retro_main_L10_while463_S2 = 1347;
  localparam retro_main_L10_while463_S3 = 1348;
  localparam retro_main_L10_ifelse566_S0 = 1349;
  localparam retro_main_L11_while470_S0 = 1350;
  localparam retro_main_L11_while470_S1 = 1351;
  localparam retro_main_L11_while470_S2 = 1352;
  localparam retro_main_L11_while470_S3 = 1353;
  localparam retro_main_L11_ifelse565_S0 = 1354;
  localparam retro_main_L12_while475_S0 = 1355;
  localparam retro_main_L12_while475_S1 = 1356;
  localparam retro_main_L12_while475_S2 = 1357;
  localparam retro_main_L12_while475_S3 = 1358;
  localparam retro_main_L12_ifelse564_S0 = 1359;
  localparam retro_main_L13_while480_S0 = 1360;
  localparam retro_main_L13_while480_S1 = 1361;
  localparam retro_main_L13_while480_S2 = 1362;
  localparam retro_main_L13_while480_S3 = 1363;
  localparam retro_main_L13_ifelse563_S0 = 1364;
  localparam retro_main_L14_while487_S0 = 1365;
  localparam retro_main_L14_while487_S1 = 1366;
  localparam retro_main_L14_while487_S2 = 1367;
  localparam retro_main_L14_while487_S3 = 1368;
  localparam retro_main_L14_ifelse562_S0 = 1369;
  localparam retro_main_L15_while492_S0 = 1370;
  localparam retro_main_L15_while492_S1 = 1371;
  localparam retro_main_L15_while492_S2 = 1372;
  localparam retro_main_L15_while492_S3 = 1373;
  localparam retro_main_L15_ifelse561_S0 = 1374;
  localparam retro_main_L16_while497_S0 = 1375;
  localparam retro_main_L16_while497_S1 = 1376;
  localparam retro_main_L16_while497_S2 = 1377;
  localparam retro_main_L16_while497_S3 = 1378;
  localparam retro_main_L16_ifelse560_S0 = 1379;
  localparam retro_main_L17_while505_S0 = 1380;
  localparam retro_main_L17_while505_S1 = 1381;
  localparam retro_main_L17_while505_S2 = 1382;
  localparam retro_main_L17_while505_S3 = 1383;
  localparam retro_main_L17_ifelse559_S0 = 1384;
  localparam retro_main_L18_while510_S0 = 1385;
  localparam retro_main_L18_while510_S1 = 1386;
  localparam retro_main_L18_while510_S2 = 1387;
  localparam retro_main_L18_while510_S3 = 1388;
  localparam retro_main_L18_ifelse558_S0 = 1389;
  localparam retro_main_L19_while515_S0 = 1390;
  localparam retro_main_L19_while515_S1 = 1391;
  localparam retro_main_L19_while515_S2 = 1392;
  localparam retro_main_L19_while515_S3 = 1393;
  localparam retro_main_L19_ifelse557_S0 = 1394;
  localparam retro_main_L20_fortest393_S0 = 1395;
  localparam retro_main_L20_forbody394_S0 = 1396;
  localparam retro_main_L20_ifelse416_S0 = 1397;
  localparam retro_main_L20_ifelse416_S1 = 1398;
  localparam retro_main_L21_fortest399_S0 = 1399;
  localparam retro_main_L21_forbody400_S0 = 1400;
  localparam retro_main_L21_ifelse414_S0 = 1401;
  localparam retro_main_L21_ifelse414_S1 = 1402;
  localparam retro_main_L22_fortest404_S0 = 1403;
  localparam retro_main_L22_forbody405_S0 = 1404;
  localparam retro_main_L22_forbody405_S1 = 1405;
  
  //signals: 
  reg        [31:0] array995_inl49 [0:1];
  reg        [31:0] array998 [0:11];
  wire c1084_inl51;
  wire c1085_inl51;
  wire c1086_inl51;
  wire c1087_inl51;
  wire c1088_inl51;
  wire c1089_inl51;
  wire c1090_inl51;
  wire c1091_inl51;
  wire c1092_inl51;
  wire c1093_inl51;
  wire c1094_inl51;
  wire c1095_inl51;
  wire c1096_inl51;
  wire c1097_inl51;
  wire c1098_inl51;
  wire c1099_inl51;
  wire c1100_inl51;
  wire c1101_inl51;
  wire c1102_inl51;
  wire c1103_inl51;
  wire c1104_inl51;
  wire c1105_inl51;
  wire c1106;
  wire c1107;
  wire c1108;
  wire c1109;
  wire c1110;
  wire c1111;
  wire c1112;
  wire c1113;
  wire c1114;
  wire c1115;
  wire c1116;
  wire c1117;
  wire c1118;
  wire c1119;
  wire c1120;
  wire c1121;
  wire c1122;
  wire c1123;
  wire c1124;
  wire c1125;
  wire c1126;
  wire c1127;
  wire c1128;
  wire c1129;
  wire c1130;
  wire c1131;
  wire c1132;
  wire c1133;
  wire c1134;
  wire c1135;
  wire c1136;
  wire c2157;
  wire c2158;
  wire c2159;
  wire c2160;
  wire c2161;
  wire c2162;
  wire c2163;
  wire c2164;
  wire c2165;
  wire c2166;
  wire c2167;
  wire c2168;
  wire c2169;
  wire c2170;
  wire c2171;
  wire c2172;
  wire c2173;
  wire c2174;
  wire c2175;
  wire c2176;
  wire c2177;
  wire c2178;
  wire c2179;
  wire c2180;
  wire c2181;
  wire c2182;
  wire c2183;
  wire c2184;
  wire c2185;
  wire c2186;
  wire c2187;
  wire c2188;
  wire c2212;
  wire c2217;
  wire c2235;
  wire c2243;
  wire c2246;
  wire c2247;
  wire c2256;
  wire c2257;
  wire c2275;
  wire c2277;
  wire c2278;
  wire c2279;
  wire c2280;
  wire c2282;
  wire c2283;
  wire c2284;
  wire c2285;
  wire c2286;
  wire c2287;
  wire c2288;
  wire c2289;
  wire c2290;
  wire c2291;
  wire c2292;
  wire c2293;
  wire c2294;
  wire c2295;
  wire c2296;
  wire c2297;
  wire c2298;
  wire c2299;
  wire c2300;
  wire c2301;
  wire c2310;
  wire c2311;
  wire c2312;
  wire c2313;
  wire c2314;
  wire c2315;
  wire c2316;
  wire c2317;
  wire c2318;
  wire c2319;
  wire c2320;
  wire c2322;
  wire c2323;
  wire c2324;
  wire c2325;
  wire c2326;
  wire c2327;
  wire c2328;
  wire c2329;
  wire c2330;
  wire c2331;
  wire c2332;
  wire c2333;
  wire c2334;
  wire c2335;
  wire c2336;
  wire c2337;
  wire c2338;
  wire c2339;
  wire c2340;
  wire c2341;
  wire c2342;
  wire c2343;
  wire c2344;
  wire c2345;
  wire c2346;
  wire c2347;
  wire c2348;
  wire c2349;
  wire c2350;
  wire c2351;
  wire c2352;
  wire c2353;
  wire c2354;
  wire c2355;
  wire c2356;
  wire c2357;
  wire c2358;
  wire c2359;
  wire c2360;
  wire c2361;
  wire c2856;
  wire c2857;
  wire c2858;
  wire c2859;
  wire c2860;
  wire c2861;
  wire c2862;
  wire c2863;
  wire c2864;
  wire c2865;
  wire c2866;
  wire c2867;
  wire c2868;
  wire c2869;
  wire c2870;
  wire c2871;
  wire c2872;
  wire c2873;
  wire c2874;
  wire c2875;
  wire c2876;
  wire c2877;
  wire c2878;
  wire c2879;
  wire c2880;
  wire c2881;
  wire c2882;
  wire c2883;
  wire c2884;
  wire c2885;
  wire c2886;
  wire c2887;
  wire c2888;
  wire c2889;
  wire c2890;
  wire c2891;
  wire c2892;
  wire c2893;
  wire c2894;
  wire c2895;
  wire c2896;
  wire c2897;
  wire c2898;
  wire c2899;
  wire c2900;
  wire c2901;
  wire c2902;
  wire c2903;
  wire c2904;
  wire c2905;
  wire c2906;
  wire c2907;
  wire c2908;
  wire c2909;
  wire c2910;
  wire c2911;
  wire c2912;
  wire c2913;
  wire c2914;
  wire c2915;
  wire c2916;
  wire c2917;
  wire c2918;
  wire c2919;
  wire c2920;
  wire c2921;
  wire c2922;
  wire c2923;
  wire c2924;
  wire c2925;
  wire c2926;
  wire c2927;
  wire c2928;
  wire c2929;
  wire c2930;
  wire c2931;
  wire c2932;
  wire c2933;
  wire c2934;
  wire c2935;
  wire c2936;
  wire c2937;
  wire c2938;
  wire c2939;
  wire c2940;
  wire c2941;
  wire c2942;
  wire c2943;
  wire c2944;
  wire c2945;
  wire c2946;
  wire c2947;
  wire c2948;
  wire c2949;
  wire c2950;
  wire c2951;
  wire c2952;
  wire c2953;
  wire c2954;
  wire c2955;
  wire c2956;
  wire c2957;
  wire c2958;
  wire c2959;
  wire c2960;
  wire c2961;
  wire c2962;
  wire c2963;
  wire c2964;
  wire c2965;
  wire c2966;
  wire c2967;
  wire c2968;
  wire c2969;
  wire c2970;
  wire c2971;
  wire c848_inl51;
  wire c851_inl51;
  wire c853_inl51;
  wire c854_inl51;
  wire c855_inl51;
  wire c856_inl51;
  wire c857_inl51;
  wire c860_inl51;
  wire c862_inl51;
  wire c864_inl51;
  wire c866_inl51;
  wire c868_inl51;
  wire c870_inl51;
  wire c872_inl51;
  wire c874_inl51;
  wire c876_inl51;
  wire c878_inl51;
  wire c880_inl51;
  wire c882_inl51;
  wire c884_inl51;
  wire c886_inl51;
  wire c888_inl51;
  wire c890_inl51;
  wire c892_inl51;
  wire c894_inl51;
  wire c896_inl51;
  wire c898_inl51;
  wire c900_inl51;
  wire c902_inl51;
  wire c904_inl51;
  wire c906_inl51;
  wire c908_inl51;
  wire c910_inl51;
  wire c914;
  wire c915;
  wire c916;
  wire c917;
  wire c918;
  wire c919;
  wire c920;
  wire c921;
  wire c922;
  wire c923;
  wire c924;
  wire c925;
  wire c926;
  wire c927;
  wire c928;
  wire c929;
  wire c930;
  wire c931;
  wire c932;
  wire c933;
  wire c934;
  wire c935;
  wire c936;
  wire c937;
  wire c938;
  wire c939;
  wire c940;
  wire c941;
  wire c942;
  wire c943;
  wire c944;
  wire c945;
  wire c946;
  wire c950;
  wire c951;
  wire c952;
  wire c955;
  wire c957;
  wire c959;
  wire c961;
  wire c964;
  wire c967;
  wire c973_inl49;
  wire c974_inl49;
  wire c975_inl49;
  wire c977_inl49;
  wire c985_inl2_inl1_inl51;
  wire c985_inl2_inl5_inl51;
  wire c985_inl2_inl6_inl51;
  wire c985_inl2_inl7_inl51;
  wire c985_inl2_inl8_inl51;
  wire c985_inl2_inl9_inl51;
  wire c985_inl3_inl1_inl51;
  wire c985_inl3_inl5_inl51;
  wire c985_inl3_inl6_inl51;
  wire c985_inl3_inl7_inl51;
  wire c985_inl3_inl8_inl51;
  wire c985_inl3_inl9_inl51;
  wire c986_inl1_inl49;
  wire c986_inl2_inl49;
  wire c988_inl1_inl49;
  wire c988_inl2_inl49;
  wire c994_inl1_inl1_inl51;
  wire c994_inl1_inl5_inl51;
  wire c994_inl1_inl6_inl51;
  wire c994_inl1_inl7_inl51;
  wire c994_inl1_inl8_inl51;
  wire c994_inl1_inl9_inl51;
  wire        [31:0] cmd_reply_inl1_inl1_inl51;
  wire        [31:0] cmd_reply_inl1_inl5_inl51;
  wire        [31:0] cmd_reply_inl1_inl6_inl51;
  wire        [31:0] cmd_reply_inl1_inl7_inl51;
  wire        [31:0] cmd_reply_inl1_inl8_inl51;
  wire        [31:0] cmd_reply_inl1_inl9_inl51;
  wire        [31:0] cmd_reply_inl2_inl1_inl51;
  wire        [31:0] cmd_reply_inl2_inl5_inl51;
  wire        [31:0] cmd_reply_inl2_inl6_inl51;
  wire        [31:0] cmd_reply_inl2_inl7_inl51;
  wire        [31:0] cmd_reply_inl2_inl8_inl51;
  wire        [31:0] cmd_reply_inl2_inl9_inl51;
  wire        [31:0] cmd_reply_inl3_inl1_inl51;
  wire        [31:0] cmd_reply_inl3_inl5_inl51;
  wire        [31:0] cmd_reply_inl3_inl6_inl51;
  wire        [31:0] cmd_reply_inl3_inl7_inl51;
  wire        [31:0] cmd_reply_inl3_inl8_inl51;
  wire        [31:0] cmd_reply_inl3_inl9_inl51;
  wire        [31:0] retro_divmod_result492 [0:1];
  wire        [31:0] t987_inl1_inl49;
  wire        [31:0] t987_inl2_inl49;
  wire        [31:0] t993_inl1_inl1_inl51;
  wire        [31:0] t993_inl1_inl5_inl51;
  wire        [31:0] t993_inl1_inl6_inl51;
  wire        [31:0] t993_inl1_inl7_inl51;
  wire        [31:0] t993_inl1_inl8_inl51;
  wire        [31:0] t993_inl1_inl9_inl51;
  wire        [31:0] test_bit_inl1_inl494;
  wire        [31:0] test_bit_inl2_inl494;
  wire        [31:0] x_inl1_inl49;
  wire        [31:0] x_inl2_inl49;
  reg        [10:0] retro_main_state;
  reg        [31:0] test_bit_inl1_inl493;
  reg        [31:0] test_bit_inl2_inl493;
  wire signed [31:0] abs_a_inl492;
  wire signed [31:0] abs_a_inl494;
  wire signed [31:0] abs_a_inl495;
  wire signed [31:0] abs_a_inl496;
  wire signed [31:0] abs_a_inl497;
  wire signed [31:0] abs_b_inl492;
  wire signed [31:0] abs_b_inl493;
  wire signed [31:0] abs_b_inl495;
  wire signed [31:0] address0_pos3;
  wire signed [31:0] address0_pos4;
  wire signed [31:0] address0_pos5;
  wire signed [31:0] address0_pos6;
  wire signed [31:0] address0_pos7;
  wire signed [31:0] address0_pos8;
  wire signed [31:0] address0_second8;
  wire signed [31:0] address0_top8;
  wire signed [31:0] c_bit_inl494;
  wire signed [31:0] c_bit_inl495;
  wire signed [31:0] c_bit_inl496;
  wire signed [31:0] c_bit_inl497;
  wire signed [31:0] c_bit_inl498;
  wire signed [31:0] c_bit_inl499;
  wire signed [31:0] find_zero_len_result2_inl494;
  wire signed [31:0] i_inl1_inl494;
  wire signed [31:0] i_inl2_inl494;
  wire signed [31:0] i_inl494;
  wire signed [31:0] ip10;
  wire signed [31:0] ip11;
  wire signed [31:0] ip12;
  wire signed [31:0] ip13;
  wire signed [31:0] ip14;
  wire signed [31:0] ip15;
  wire signed [31:0] ip16;
  wire signed [31:0] ip17;
  wire signed [31:0] ip20;
  wire signed [31:0] ip21;
  wire signed [31:0] ip22;
  wire signed [31:0] ip3;
  wire signed [31:0] ip4;
  wire signed [31:0] ip5;
  wire signed [31:0] ip6;
  wire signed [31:0] ip7;
  wire signed [31:0] ip8;
  wire signed [31:0] ip_inl514;
  wire signed [31:0] n_inl1_inl494;
  wire signed [31:0] n_inl2_inl494;
  wire signed [31:0] stack0_pos10;
  wire signed [31:0] stack0_pos11;
  wire signed [31:0] stack0_pos12;
  wire signed [31:0] stack0_pos13;
  wire signed [31:0] stack0_pos14;
  wire signed [31:0] stack0_pos15;
  wire signed [31:0] stack0_pos16;
  wire signed [31:0] stack0_pos17;
  wire signed [31:0] stack0_pos18;
  wire signed [31:0] stack0_pos19;
  wire signed [31:0] stack0_pos20;
  wire signed [31:0] stack0_pos21;
  wire signed [31:0] stack0_pos22;
  wire signed [31:0] stack0_pos23;
  wire signed [31:0] stack0_pos24;
  wire signed [31:0] stack0_pos25;
  wire signed [31:0] stack0_pos26;
  wire signed [31:0] stack0_pos27;
  wire signed [31:0] stack0_pos28;
  wire signed [31:0] stack0_pos29;
  wire signed [31:0] stack0_pos30;
  wire signed [31:0] stack0_pos31;
  wire signed [31:0] stack0_pos32;
  wire signed [31:0] stack0_pos33;
  wire signed [31:0] stack0_pos34;
  wire signed [31:0] stack0_pos35;
  wire signed [31:0] stack0_pos3;
  wire signed [31:0] stack0_pos4;
  wire signed [31:0] stack0_pos5;
  wire signed [31:0] stack0_pos6;
  wire signed [31:0] stack0_pos7;
  wire signed [31:0] stack0_pos8;
  wire signed [31:0] stack0_pos9;
  wire signed [31:0] stack0_second23;
  wire signed [31:0] stack0_second35;
  wire signed [31:0] stack0_second36;
  wire signed [31:0] stack0_second37;
  wire signed [31:0] stack0_top23;
  wire signed [31:0] stack0_top25;
  wire signed [31:0] stack0_top27;
  wire signed [31:0] stack0_top28;
  wire signed [31:0] stack0_top30;
  wire signed [31:0] stack0_top32;
  wire signed [31:0] stack0_top34;
  wire signed [31:0] stack0_top36;
  wire signed [31:0] stack0_top38;
  wire signed [31:0] stack0_top40;
  wire signed [31:0] stack0_top41;
  wire signed [31:0] stack0_top49;
  wire signed [31:0] stack0_top50;
  wire signed [31:0] stack0_top9;
  wire signed [31:0] t2660;
  wire signed [31:0] t2670;
  wire signed [31:0] t2680;
  wire signed [31:0] t2690;
  wire signed [31:0] t486_inl49;
  wire signed [31:0] t843_inl3;
  wire signed [31:0] t843_inl4;
  wire signed [31:0] t843_inl5;
  wire signed [31:0] t843_inl6;
  wire signed [31:0] t843_inl7;
  wire signed [31:0] t846_inl10;
  wire signed [31:0] t846_inl11;
  wire signed [31:0] t846_inl12;
  wire signed [31:0] t846_inl13;
  wire signed [31:0] t846_inl14;
  wire signed [31:0] t846_inl15;
  wire signed [31:0] t846_inl16;
  wire signed [31:0] t846_inl17;
  wire signed [31:0] t846_inl18;
  wire signed [31:0] t846_inl19;
  wire signed [31:0] t846_inl20;
  wire signed [31:0] t846_inl21;
  wire signed [31:0] t846_inl22;
  wire signed [31:0] t846_inl23;
  wire signed [31:0] t846_inl24;
  wire signed [31:0] t846_inl25;
  wire signed [31:0] t846_inl26;
  wire signed [31:0] t846_inl27;
  wire signed [31:0] t846_inl28;
  wire signed [31:0] t846_inl29;
  wire signed [31:0] t846_inl2_inl51;
  wire signed [31:0] t846_inl30;
  wire signed [31:0] t846_inl31;
  wire signed [31:0] t846_inl32;
  wire signed [31:0] t846_inl33;
  wire signed [31:0] t846_inl34;
  wire signed [31:0] t846_inl3_inl51;
  wire signed [31:0] t846_inl4_inl51;
  wire signed [31:0] t846_inl8;
  wire signed [31:0] t846_inl9;
  wire signed [31:0] t969_inl49;
  wire signed [31:0] t970_inl49;
  wire signed [31:0] t971_inl49;
  wire signed [31:0] t972_inl49;
  wire signed [31:0] t976_inl49;
  reg signed [31:0] a6;
  reg signed [31:0] abs_a_inl493;
  reg signed [31:0] abs_b_inl494;
  reg signed [31:0] address0_pos2;
  reg signed [31:0] address0_second2;
  reg signed [31:0] address0_second4;
  reg signed [31:0] address0_second5;
  reg signed [31:0] address0_second6;
  reg signed [31:0] address0_top2;
  reg signed [31:0] b6;
  reg signed [31:0] c_bit_inl493;
  reg signed [31:0] char_c_inl1_inl51;
  reg signed [31:0] i_inl1_inl493;
  reg signed [31:0] i_inl2_inl493;
  reg signed [31:0] i_inl493;
  reg signed [31:0] ip2;
  reg signed [31:0] n_inl1_inl493;
  reg signed [31:0] n_inl2_inl493;
  reg signed [31:0] opcode3;
  reg signed [31:0] stack0_pos2;
  reg signed [31:0] stack0_second10;
  reg signed [31:0] stack0_second11;
  reg signed [31:0] stack0_second12;
  reg signed [31:0] stack0_second13;
  reg signed [31:0] stack0_second14;
  reg signed [31:0] stack0_second15;
  reg signed [31:0] stack0_second16;
  reg signed [31:0] stack0_second17;
  reg signed [31:0] stack0_second18;
  reg signed [31:0] stack0_second19;
  reg signed [31:0] stack0_second20;
  reg signed [31:0] stack0_second21;
  reg signed [31:0] stack0_second22;
  reg signed [31:0] stack0_second24;
  reg signed [31:0] stack0_second25;
  reg signed [31:0] stack0_second26;
  reg signed [31:0] stack0_second27;
  reg signed [31:0] stack0_second28;
  reg signed [31:0] stack0_second29;
  reg signed [31:0] stack0_second2;
  reg signed [31:0] stack0_second30;
  reg signed [31:0] stack0_second31;
  reg signed [31:0] stack0_second32;
  reg signed [31:0] stack0_second33;
  reg signed [31:0] stack0_second34;
  reg signed [31:0] stack0_second5;
  reg signed [31:0] stack0_second7;
  reg signed [31:0] stack0_second9;
  reg signed [31:0] stack0_top19;
  reg signed [31:0] stack0_top2;
  reg signed [31:0] stack0_top42;
  reg signed [31:0] t11;
  reg signed [31:0] t847_inl51;
  reg signed [31:0] t850_inl51;
  reg signed [31:0] t852_inl51;
  reg signed [31:0] t859_inl51;
  reg signed [31:0] t861_inl51;
  reg signed [31:0] t863_inl51;
  reg signed [31:0] t865_inl51;
  reg signed [31:0] t867_inl51;
  reg signed [31:0] t869_inl51;
  reg signed [31:0] t871_inl51;
  reg signed [31:0] t873_inl51;
  reg signed [31:0] t875_inl51;
  reg signed [31:0] t877_inl51;
  reg signed [31:0] t879_inl51;
  reg signed [31:0] t881_inl51;
  reg signed [31:0] t883_inl51;
  reg signed [31:0] t885_inl51;
  reg signed [31:0] t887_inl51;
  reg signed [31:0] t889_inl51;
  reg signed [31:0] t891_inl51;
  reg signed [31:0] t893_inl51;
  reg signed [31:0] t895_inl51;
  reg signed [31:0] t897_inl51;
  reg signed [31:0] t899_inl51;
  reg signed [31:0] t901_inl51;
  reg signed [31:0] t903_inl51;
  reg signed [31:0] t905_inl51;
  reg signed [31:0] t907_inl51;
  reg signed [31:0] t909_inl51;
  reg signed [31:0] t947;
  reg signed [31:0] t953;
  reg signed [31:0] t954;
  reg signed [31:0] t956;
  reg signed [31:0] t958;
  reg signed [31:0] t960;
  reg signed [31:0] t962;
  reg signed [31:0] t966;
  reg signed [31:0] t968;
  reg signed [31:0] t983_inl2_inl1_inl51;
  reg signed [31:0] t983_inl2_inl5_inl51;
  reg signed [31:0] t983_inl2_inl6_inl51;
  reg signed [31:0] t983_inl2_inl7_inl51;
  reg signed [31:0] t983_inl2_inl8_inl51;
  reg signed [31:0] t983_inl2_inl9_inl51;
  reg signed [31:0] t983_inl3_inl1_inl51;
  reg signed [31:0] t983_inl3_inl5_inl51;
  reg signed [31:0] t983_inl3_inl6_inl51;
  reg signed [31:0] t983_inl3_inl7_inl51;
  reg signed [31:0] t983_inl3_inl8_inl51;
  reg signed [31:0] t983_inl3_inl9_inl51;
  reg signed [31:0] t992_inl1_inl1_inl51;
  reg signed [31:0] t992_inl1_inl5_inl51;
  reg signed [31:0] t992_inl1_inl6_inl51;
  reg signed [31:0] t992_inl1_inl7_inl51;
  reg signed [31:0] t992_inl1_inl8_inl51;
  reg signed [31:0] t992_inl1_inl9_inl51;
  //signals: _address
  wire        [10:0] _address_len;
  wire        [31:0] _address_q;
  reg        [10:0] _address_addr;
  reg        [31:0] _address_d;
  reg _address_req;
  reg _address_we;
  //signals: _stack
  wire        [7:0] _stack_len;
  wire        [31:0] _stack_q;
  reg        [7:0] _stack_addr;
  reg        [31:0] _stack_d;
  reg _stack_req;
  reg _stack_we;
  //signals: io_ports
  wire        [4:0] io_ports_len;
  wire        [31:0] io_ports_q;
  reg        [4:0] io_ports_addr;
  reg        [31:0] io_ports_d;
  reg io_ports_req;
  reg io_ports_we;
  //signals: memory
  wire        [14:0] memory_len;
  wire        [31:0] memory_q;
  reg        [14:0] memory_addr;
  reg        [31:0] memory_d;
  reg memory_req;
  reg memory_we;
  //signals: ram
  wire        [7:0] array996_ram_addr;
  wire        [31:0] array996_ram_d;
  wire        [7:0] array996_ram_len;
  wire        [31:0] array996_ram_q;
  wire array996_ram_we;
  wire        [10:0] array997_ram_addr;
  wire        [31:0] array997_ram_d;
  wire        [10:0] array997_ram_len;
  wire        [31:0] array997_ram_q;
  wire array997_ram_we;
  //combinations: 
  assign abs_a_inl492 = (stack0_second2 & 2147483647);
  assign abs_a_inl494 = (abs_a_inl493 | 2147483648);
  assign abs_a_inl495 = c2294 ? abs_a_inl494 : ((c2286 || c2284) && !c975_inl49) ? abs_a_inl493 : 'bz;
  assign abs_a_inl496 = (abs_a_inl493 - abs_b_inl494);
  assign abs_a_inl497 = c2292 ? abs_a_inl496 : c2293 ? abs_a_inl493 : 'bz;
  assign abs_b_inl492 = (stack0_top2 & 2147483647);
  assign abs_b_inl493 = (abs_b_inl492 << find_zero_len_result2_inl494);
  assign abs_b_inl495 = (abs_b_inl494 >>> 1);
  assign address0_pos3 = (address0_pos2 + 1);
  assign address0_pos4 = (address0_pos2 - 1);
  assign address0_pos5 = (address0_pos2 - 1);
  assign address0_pos6 = (address0_pos2 - 1);
  assign address0_pos7 = (address0_pos2 + 1);
  assign address0_pos8 = (c2157 && c916) ? address0_pos2 : c2159 ? address0_pos2 : c2160 ? address0_pos2 : c2161 ? address0_pos2 : c2162 ? address0_pos2 : c2163 ? address0_pos3 : c2164 ? address0_pos4 : c2246 ? address0_pos2 : c2247 ? address0_pos2 : c2166 ? address0_pos2 : c2167 ? address0_pos5 : c2168 ? address0_pos2 : c2169 ? address0_pos2 : c2170 ? address0_pos2 : c2171 ? address0_pos2 : c2172 ? address0_pos2 : c2173 ? address0_pos2 : c2174 ? address0_pos2 : c2175 ? address0_pos2 : c2176 ? address0_pos2 : (c2286 || c2284) ? address0_pos2 : c2178 ? address0_pos2 : c2179 ? address0_pos2 : c2180 ? address0_pos2 : c2181 ? address0_pos2 : c2182 ? address0_pos2 : c2212 ? address0_pos6 : (c2183 && !c964) ? address0_pos2 : c2184 ? address0_pos2 : c2185 ? address0_pos2 : c2186 ? address0_pos2 : c2187 ? address0_pos2 : (c2361 || c2360) ? address0_pos2 : (c2188 && !c967) ? address0_pos2 : (c2157 && c1136) ? address0_pos2 : c2158 ? address0_pos7 : 'bz;
  assign address0_second8 = (c2157 && c916) ? address0_second2 : c2159 ? address0_second2 : c2160 ? address0_second2 : c2161 ? address0_second2 : c2162 ? address0_second2 : c2163 ? address0_top2 : c2164 ? address0_second4 : c2246 ? address0_second2 : c2247 ? address0_second2 : c2166 ? address0_second2 : c2167 ? address0_second5 : c2168 ? address0_second2 : c2169 ? address0_second2 : c2170 ? address0_second2 : c2171 ? address0_second2 : c2172 ? address0_second2 : c2173 ? address0_second2 : c2174 ? address0_second2 : c2175 ? address0_second2 : c2176 ? address0_second2 : (c2286 || c2284) ? address0_second2 : c2178 ? address0_second2 : c2179 ? address0_second2 : c2180 ? address0_second2 : c2181 ? address0_second2 : c2182 ? address0_second2 : c2212 ? address0_second6 : (c2183 && !c964) ? address0_second2 : c2184 ? address0_second2 : c2185 ? address0_second2 : c2186 ? address0_second2 : c2187 ? address0_second2 : (c2361 || c2360) ? address0_second2 : (c2188 && !c967) ? address0_second2 : (c2157 && c1136) ? address0_second2 : c2158 ? address0_top2 : 'bz;
  assign address0_top8 = (c2157 && c916) ? address0_top2 : c2159 ? address0_top2 : c2160 ? address0_top2 : c2161 ? address0_top2 : c2162 ? address0_top2 : c2163 ? stack0_top2 : c2164 ? address0_second2 : c2246 ? address0_top2 : c2247 ? address0_top2 : c2166 ? address0_top2 : c2167 ? address0_second2 : c2168 ? address0_top2 : c2169 ? address0_top2 : c2170 ? address0_top2 : c2171 ? address0_top2 : c2172 ? address0_top2 : c2173 ? address0_top2 : c2174 ? address0_top2 : c2175 ? address0_top2 : c2176 ? address0_top2 : (c2286 || c2284) ? address0_top2 : c2178 ? address0_top2 : c2179 ? address0_top2 : c2180 ? address0_top2 : c2181 ? address0_top2 : c2182 ? address0_top2 : c2212 ? address0_second2 : (c2183 && !c964) ? address0_top2 : c2184 ? address0_top2 : c2185 ? address0_top2 : c2186 ? address0_top2 : c2187 ? address0_top2 : (c2361 || c2360) ? address0_top2 : (c2188 && !c967) ? address0_top2 : (c2157 && c1136) ? address0_top2 : c2158 ? ip2 : 'bz;
  assign c1084_inl51 = (!c864_inl51 && c866_inl51);
  assign c1085_inl51 = ((!c864_inl51 && !c866_inl51) && c868_inl51);
  assign c1086_inl51 = (((!c864_inl51 && !c866_inl51) && !c868_inl51) && c870_inl51);
  assign c1087_inl51 = ((((!c864_inl51 && !c866_inl51) && !c868_inl51) && !c870_inl51) && c872_inl51);
  assign c1088_inl51 = (((((!c864_inl51 && !c866_inl51) && !c868_inl51) && !c870_inl51) && !c872_inl51) && c874_inl51);
  assign c1089_inl51 = ((((((!c864_inl51 && !c866_inl51) && !c868_inl51) && !c870_inl51) && !c872_inl51) && !c874_inl51) && c876_inl51);
  assign c1090_inl51 = ((((((!c864_inl51 && !c866_inl51) && !c868_inl51) && !c870_inl51) && !c872_inl51) && !c874_inl51) && !c876_inl51);
  assign c1091_inl51 = (!c880_inl51 && c882_inl51);
  assign c1092_inl51 = ((!c880_inl51 && !c882_inl51) && c884_inl51);
  assign c1093_inl51 = (((!c880_inl51 && !c882_inl51) && !c884_inl51) && c886_inl51);
  assign c1094_inl51 = ((((!c880_inl51 && !c882_inl51) && !c884_inl51) && !c886_inl51) && c888_inl51);
  assign c1095_inl51 = (((((!c880_inl51 && !c882_inl51) && !c884_inl51) && !c886_inl51) && !c888_inl51) && c890_inl51);
  assign c1096_inl51 = ((((((!c880_inl51 && !c882_inl51) && !c884_inl51) && !c886_inl51) && !c888_inl51) && !c890_inl51) && c892_inl51);
  assign c1097_inl51 = (((((((!c880_inl51 && !c882_inl51) && !c884_inl51) && !c886_inl51) && !c888_inl51) && !c890_inl51) && !c892_inl51) && c894_inl51);
  assign c1098_inl51 = ((((((((!c880_inl51 && !c882_inl51) && !c884_inl51) && !c886_inl51) && !c888_inl51) && !c890_inl51) && !c892_inl51) && !c894_inl51) && c896_inl51);
  assign c1099_inl51 = (((((((((!c880_inl51 && !c882_inl51) && !c884_inl51) && !c886_inl51) && !c888_inl51) && !c890_inl51) && !c892_inl51) && !c894_inl51) && !c896_inl51) && c898_inl51);
  assign c1100_inl51 = ((((((((((!c880_inl51 && !c882_inl51) && !c884_inl51) && !c886_inl51) && !c888_inl51) && !c890_inl51) && !c892_inl51) && !c894_inl51) && !c896_inl51) && !c898_inl51) && c900_inl51);
  assign c1101_inl51 = (((((((((((!c880_inl51 && !c882_inl51) && !c884_inl51) && !c886_inl51) && !c888_inl51) && !c890_inl51) && !c892_inl51) && !c894_inl51) && !c896_inl51) && !c898_inl51) && !c900_inl51) && c902_inl51);
  assign c1102_inl51 = ((((((((((((!c880_inl51 && !c882_inl51) && !c884_inl51) && !c886_inl51) && !c888_inl51) && !c890_inl51) && !c892_inl51) && !c894_inl51) && !c896_inl51) && !c898_inl51) && !c900_inl51) && !c902_inl51) && c904_inl51);
  assign c1103_inl51 = (((((((((((((!c880_inl51 && !c882_inl51) && !c884_inl51) && !c886_inl51) && !c888_inl51) && !c890_inl51) && !c892_inl51) && !c894_inl51) && !c896_inl51) && !c898_inl51) && !c900_inl51) && !c902_inl51) && !c904_inl51) && c906_inl51);
  assign c1104_inl51 = ((((((((((((((!c880_inl51 && !c882_inl51) && !c884_inl51) && !c886_inl51) && !c888_inl51) && !c890_inl51) && !c892_inl51) && !c894_inl51) && !c896_inl51) && !c898_inl51) && !c900_inl51) && !c902_inl51) && !c904_inl51) && !c906_inl51) && c908_inl51);
  assign c1105_inl51 = ((((((((((((((!c880_inl51 && !c882_inl51) && !c884_inl51) && !c886_inl51) && !c888_inl51) && !c890_inl51) && !c892_inl51) && !c894_inl51) && !c896_inl51) && !c898_inl51) && !c900_inl51) && !c902_inl51) && !c904_inl51) && !c906_inl51) && !c908_inl51);
  assign c1106 = (!c916 && c917);
  assign c1107 = ((!c916 && !c917) && c918);
  assign c1108 = (((!c916 && !c917) && !c918) && c919);
  assign c1109 = ((((!c916 && !c917) && !c918) && !c919) && c920);
  assign c1110 = (((((!c916 && !c917) && !c918) && !c919) && !c920) && c921);
  assign c1111 = ((((((!c916 && !c917) && !c918) && !c919) && !c920) && !c921) && c922);
  assign c1112 = (((((((!c916 && !c917) && !c918) && !c919) && !c920) && !c921) && !c922) && c923);
  assign c1113 = ((((((((!c916 && !c917) && !c918) && !c919) && !c920) && !c921) && !c922) && !c923) && c924);
  assign c1114 = (((((((((!c916 && !c917) && !c918) && !c919) && !c920) && !c921) && !c922) && !c923) && !c924) && c925);
  assign c1115 = ((((((((((!c916 && !c917) && !c918) && !c919) && !c920) && !c921) && !c922) && !c923) && !c924) && !c925) && c926);
  assign c1116 = (((((((((((!c916 && !c917) && !c918) && !c919) && !c920) && !c921) && !c922) && !c923) && !c924) && !c925) && !c926) && c927);
  assign c1117 = ((((((((((((!c916 && !c917) && !c918) && !c919) && !c920) && !c921) && !c922) && !c923) && !c924) && !c925) && !c926) && !c927) && c928);
  assign c1118 = (((((((((((((!c916 && !c917) && !c918) && !c919) && !c920) && !c921) && !c922) && !c923) && !c924) && !c925) && !c926) && !c927) && !c928) && c929);
  assign c1119 = ((((((((((((((!c916 && !c917) && !c918) && !c919) && !c920) && !c921) && !c922) && !c923) && !c924) && !c925) && !c926) && !c927) && !c928) && !c929) && c930);
  assign c1120 = (((((((((((((((!c916 && !c917) && !c918) && !c919) && !c920) && !c921) && !c922) && !c923) && !c924) && !c925) && !c926) && !c927) && !c928) && !c929) && !c930) && c931);
  assign c1121 = ((((((((((((((((!c916 && !c917) && !c918) && !c919) && !c920) && !c921) && !c922) && !c923) && !c924) && !c925) && !c926) && !c927) && !c928) && !c929) && !c930) && !c931) && c932);
  assign c1122 = (((((((((((((((((!c916 && !c917) && !c918) && !c919) && !c920) && !c921) && !c922) && !c923) && !c924) && !c925) && !c926) && !c927) && !c928) && !c929) && !c930) && !c931) && !c932) && c933);
  assign c1123 = ((((((((((((((((((!c916 && !c917) && !c918) && !c919) && !c920) && !c921) && !c922) && !c923) && !c924) && !c925) && !c926) && !c927) && !c928) && !c929) && !c930) && !c931) && !c932) && !c933) && c934);
  assign c1124 = (((((((((((((((((((!c916 && !c917) && !c918) && !c919) && !c920) && !c921) && !c922) && !c923) && !c924) && !c925) && !c926) && !c927) && !c928) && !c929) && !c930) && !c931) && !c932) && !c933) && !c934) && c935);
  assign c1125 = ((((((((((((((((((((!c916 && !c917) && !c918) && !c919) && !c920) && !c921) && !c922) && !c923) && !c924) && !c925) && !c926) && !c927) && !c928) && !c929) && !c930) && !c931) && !c932) && !c933) && !c934) && !c935) && c936);
  assign c1126 = (((((((((((((((((((((!c916 && !c917) && !c918) && !c919) && !c920) && !c921) && !c922) && !c923) && !c924) && !c925) && !c926) && !c927) && !c928) && !c929) && !c930) && !c931) && !c932) && !c933) && !c934) && !c935) && !c936) && c937);
  assign c1127 = ((((((((((((((((((((((!c916 && !c917) && !c918) && !c919) && !c920) && !c921) && !c922) && !c923) && !c924) && !c925) && !c926) && !c927) && !c928) && !c929) && !c930) && !c931) && !c932) && !c933) && !c934) && !c935) && !c936) && !c937) && c938);
  assign c1128 = (((((((((((((((((((((((!c916 && !c917) && !c918) && !c919) && !c920) && !c921) && !c922) && !c923) && !c924) && !c925) && !c926) && !c927) && !c928) && !c929) && !c930) && !c931) && !c932) && !c933) && !c934) && !c935) && !c936) && !c937) && !c938) && c939);
  assign c1129 = ((((((((((((((((((((((((!c916 && !c917) && !c918) && !c919) && !c920) && !c921) && !c922) && !c923) && !c924) && !c925) && !c926) && !c927) && !c928) && !c929) && !c930) && !c931) && !c932) && !c933) && !c934) && !c935) && !c936) && !c937) && !c938) && !c939) && c940);
  assign c1130 = (((((((((((((((((((((((((!c916 && !c917) && !c918) && !c919) && !c920) && !c921) && !c922) && !c923) && !c924) && !c925) && !c926) && !c927) && !c928) && !c929) && !c930) && !c931) && !c932) && !c933) && !c934) && !c935) && !c936) && !c937) && !c938) && !c939) && !c940) && c941);
  assign c1131 = ((((((((((((((((((((((((((!c916 && !c917) && !c918) && !c919) && !c920) && !c921) && !c922) && !c923) && !c924) && !c925) && !c926) && !c927) && !c928) && !c929) && !c930) && !c931) && !c932) && !c933) && !c934) && !c935) && !c936) && !c937) && !c938) && !c939) && !c940) && !c941) && c942);
  assign c1132 = (((((((((((((((((((((((((((!c916 && !c917) && !c918) && !c919) && !c920) && !c921) && !c922) && !c923) && !c924) && !c925) && !c926) && !c927) && !c928) && !c929) && !c930) && !c931) && !c932) && !c933) && !c934) && !c935) && !c936) && !c937) && !c938) && !c939) && !c940) && !c941) && !c942) && c943);
  assign c1133 = ((((((((((((((((((((((((((((!c916 && !c917) && !c918) && !c919) && !c920) && !c921) && !c922) && !c923) && !c924) && !c925) && !c926) && !c927) && !c928) && !c929) && !c930) && !c931) && !c932) && !c933) && !c934) && !c935) && !c936) && !c937) && !c938) && !c939) && !c940) && !c941) && !c942) && !c943) && c944);
  assign c1134 = (((((((((((((((((((((((((((((!c916 && !c917) && !c918) && !c919) && !c920) && !c921) && !c922) && !c923) && !c924) && !c925) && !c926) && !c927) && !c928) && !c929) && !c930) && !c931) && !c932) && !c933) && !c934) && !c935) && !c936) && !c937) && !c938) && !c939) && !c940) && !c941) && !c942) && !c943) && !c944) && c945);
  assign c1135 = ((((((((((((((((((((((((((((((!c916 && !c917) && !c918) && !c919) && !c920) && !c921) && !c922) && !c923) && !c924) && !c925) && !c926) && !c927) && !c928) && !c929) && !c930) && !c931) && !c932) && !c933) && !c934) && !c935) && !c936) && !c937) && !c938) && !c939) && !c940) && !c941) && !c942) && !c943) && !c944) && !c945) && c946);
  assign c1136 = ((((((((((((((((((((((((((((((!c916 && !c917) && !c918) && !c919) && !c920) && !c921) && !c922) && !c923) && !c924) && !c925) && !c926) && !c927) && !c928) && !c929) && !c930) && !c931) && !c932) && !c933) && !c934) && !c935) && !c936) && !c937) && !c938) && !c939) && !c940) && !c941) && !c942) && !c943) && !c944) && !c945) && !c946);
  assign c2157 = (c914 && c915);
  assign c2158 = (c914 && !c915);
  assign c2159 = (c2157 && c1106);
  assign c2160 = (c2157 && c1107);
  assign c2161 = (c2157 && c1108);
  assign c2162 = (c2157 && c1109);
  assign c2163 = (c2157 && c1110);
  assign c2164 = (c2157 && c1111);
  assign c2165 = (c2157 && c1112);
  assign c2166 = (c2157 && c1113);
  assign c2167 = (c2157 && c1114);
  assign c2168 = (c2157 && c1115);
  assign c2169 = (c2157 && c1116);
  assign c2170 = (c2157 && c1117);
  assign c2171 = (c2157 && c1118);
  assign c2172 = (c2157 && c1119);
  assign c2173 = (c2157 && c1120);
  assign c2174 = (c2157 && c1121);
  assign c2175 = (c2157 && c1122);
  assign c2176 = (c2157 && c1123);
  assign c2177 = (c2157 && c1124);
  assign c2178 = (c2157 && c1125);
  assign c2179 = (c2157 && c1126);
  assign c2180 = (c2157 && c1127);
  assign c2181 = (c2157 && c1128);
  assign c2182 = (c2157 && c1129);
  assign c2183 = (c2157 && c1130);
  assign c2184 = (c2157 && c1131);
  assign c2185 = (c2157 && c1132);
  assign c2186 = (c2157 && c1133);
  assign c2187 = (c2157 && c1134);
  assign c2188 = (c2157 && c1135);
  assign c2212 = (c2183 && c964);
  assign c2217 = (c2188 && c967);
  assign c2235 = (c2177 && c986_inl1_inl49);
  assign c2243 = (c2217 && c848_inl51);
  assign c2246 = (c2165 && c952);
  assign c2247 = (c2165 && !c952);
  assign c2256 = (c2235 && c988_inl1_inl49);
  assign c2257 = (c2235 && !c988_inl1_inl49);
  assign c2275 = (c2243 && !c994_inl1_inl1_inl51);
  assign c2277 = (c2168 && c955);
  assign c2278 = (c2169 && c957);
  assign c2279 = (c2170 && c959);
  assign c2280 = (c2171 && c961);
  assign c2282 = ((c2177 || c2256) && c986_inl2_inl49);
  assign c2283 = (c2243 && !c985_inl2_inl1_inl51);
  assign c2284 = (c2282 && c988_inl2_inl49);
  assign c2285 = (c2282 && !c988_inl2_inl49);
  assign c2286 = (c2177 || c2256);
  assign c2287 = (c2243 && !c985_inl3_inl1_inl51);
  assign c2288 = (c2243 && c851_inl51);
  assign c2289 = ((c2286 || c2284) && c973_inl49);
  assign c2290 = (c2217 && !c848_inl51);
  assign c2291 = (c2243 && !c851_inl51);
  assign c2292 = (c2289 && c974_inl49);
  assign c2293 = (c2289 && !c974_inl49);
  assign c2294 = ((c2286 || c2284) && c975_inl49);
  assign c2295 = (((c2290 || c2291) || c2288) && c853_inl51);
  assign c2296 = ((c2286 || c2284) && !c975_inl49);
  assign c2297 = (c2295 && c856_inl51);
  assign c2298 = (c2295 && !c856_inl51);
  assign c2299 = ((c2296 || c2294) && c977_inl49);
  assign c2300 = (c2297 && c857_inl51);
  assign c2301 = (c2297 && !c857_inl51);
  assign c2310 = (c2300 && !c994_inl1_inl5_inl51);
  assign c2311 = (c2301 && !c994_inl1_inl8_inl51);
  assign c2312 = (c2300 && !c985_inl2_inl5_inl51);
  assign c2313 = (c2301 && !c985_inl2_inl8_inl51);
  assign c2314 = (c2300 && !c985_inl3_inl5_inl51);
  assign c2315 = (c2301 && !c985_inl3_inl8_inl51);
  assign c2316 = (c2300 && !c994_inl1_inl6_inl51);
  assign c2317 = (c2300 && !c985_inl2_inl6_inl51);
  assign c2318 = (c2300 && !c985_inl3_inl6_inl51);
  assign c2319 = (c2300 && !c994_inl1_inl7_inl51);
  assign c2320 = (c2300 && !c985_inl2_inl7_inl51);
  assign c2322 = (c2301 && c985_inl3_inl8_inl51);
  assign c2323 = (c2300 && c985_inl3_inl7_inl51);
  assign c2324 = (c2300 && !c985_inl3_inl7_inl51);
  assign c2325 = (((c2298 || c2322) || c2323) && !c994_inl1_inl9_inl51);
  assign c2326 = (((c2298 || c2322) || c2323) && !c985_inl2_inl9_inl51);
  assign c2327 = (((c2298 || c2322) || c2323) && !c985_inl3_inl9_inl51);
  assign c2328 = (((c2290 || c2291) || c2288) && !c853_inl51);
  assign c2329 = ((c2298 || c2322) || c2323);
  assign c2330 = ((c2328 || c2329) && c860_inl51);
  assign c2331 = ((c2328 || c2329) && !c860_inl51);
  assign c2332 = ((c2331 || c2330) && c862_inl51);
  assign c2333 = ((c2331 || c2330) && !c862_inl51);
  assign c2334 = ((c2333 || c2332) && c864_inl51);
  assign c2335 = ((c2333 || c2332) && c1084_inl51);
  assign c2336 = ((c2333 || c2332) && c1085_inl51);
  assign c2337 = ((c2333 || c2332) && c1086_inl51);
  assign c2338 = ((c2333 || c2332) && c1087_inl51);
  assign c2339 = ((c2333 || c2332) && c1088_inl51);
  assign c2340 = ((c2333 || c2332) && c1089_inl51);
  assign c2341 = ((c2333 || c2332) && c1090_inl51);
  assign c2342 = ((((((((c2341 || c2336) || c2334) || c2335) || c2340) || c2339) || c2338) || c2337) && c878_inl51);
  assign c2343 = ((((((((c2341 || c2336) || c2334) || c2335) || c2340) || c2339) || c2338) || c2337) && !c878_inl51);
  assign c2344 = ((c2343 || c2342) && c880_inl51);
  assign c2345 = ((c2343 || c2342) && c1091_inl51);
  assign c2346 = ((c2343 || c2342) && c1092_inl51);
  assign c2347 = ((c2343 || c2342) && c1093_inl51);
  assign c2348 = ((c2343 || c2342) && c1094_inl51);
  assign c2349 = ((c2343 || c2342) && c1095_inl51);
  assign c2350 = ((c2343 || c2342) && c1096_inl51);
  assign c2351 = ((c2343 || c2342) && c1097_inl51);
  assign c2352 = ((c2343 || c2342) && c1098_inl51);
  assign c2353 = ((c2343 || c2342) && c1099_inl51);
  assign c2354 = ((c2343 || c2342) && c1100_inl51);
  assign c2355 = ((c2343 || c2342) && c1101_inl51);
  assign c2356 = ((c2343 || c2342) && c1102_inl51);
  assign c2357 = ((c2343 || c2342) && c1103_inl51);
  assign c2358 = ((c2343 || c2342) && c1104_inl51);
  assign c2359 = ((c2343 || c2342) && c1105_inl51);
  assign c2360 = ((((((((((((((((c2359 || c2349) || c2344) || c2357) || c2348) || c2347) || c2350) || c2351) || c2356) || c2353) || c2355) || c2358) || c2354) || c2346) || c2352) || c2345) && c910_inl51);
  assign c2361 = ((((((((((((((((c2359 || c2349) || c2344) || c2357) || c2348) || c2347) || c2350) || c2351) || c2356) || c2353) || c2355) || c2358) || c2354) || c2346) || c2352) || c2345) && !c910_inl51);
  assign c2856 = (c914 && c915);
  assign c2857 = (c914 && !c915);
  assign c2858 = (c2856 && c1106);
  assign c2859 = (c2856 && c1107);
  assign c2860 = (c2856 && c1108);
  assign c2861 = (c2856 && c1109);
  assign c2862 = (c2856 && c1110);
  assign c2863 = (c2856 && c1111);
  assign c2864 = (c2856 && c1112);
  assign c2865 = (c2856 && c1113);
  assign c2866 = (c2856 && c1114);
  assign c2867 = (c2856 && c1115);
  assign c2868 = (c2856 && c1116);
  assign c2869 = (c2856 && c1117);
  assign c2870 = (c2856 && c1118);
  assign c2871 = (c2856 && c1119);
  assign c2872 = (c2856 && c1120);
  assign c2873 = (c2856 && c1121);
  assign c2874 = (c2856 && c1122);
  assign c2875 = (c2856 && c1123);
  assign c2876 = (c2856 && c1124);
  assign c2877 = (c2856 && c1125);
  assign c2878 = (c2856 && c1126);
  assign c2879 = (c2856 && c1127);
  assign c2880 = (c2856 && c1128);
  assign c2881 = (c2856 && c1129);
  assign c2882 = (c2856 && c1130);
  assign c2883 = (c2856 && c1131);
  assign c2884 = (c2856 && c1132);
  assign c2885 = (c2856 && c1133);
  assign c2886 = (c2856 && c1134);
  assign c2887 = (c2856 && c1135);
  assign c2888 = (c2864 && c952);
  assign c2889 = (c2864 && !c952);
  assign c2890 = (c2867 && c955);
  assign c2891 = (c2868 && c957);
  assign c2892 = (c2869 && c959);
  assign c2893 = (c2870 && c961);
  assign c2894 = (c2882 && c964);
  assign c2895 = (c2887 && c967);
  assign c2896 = (c2867 && !c955);
  assign c2897 = (c2868 && !c957);
  assign c2898 = (c2869 && !c959);
  assign c2899 = (c2870 && !c961);
  assign c2900 = (c2876 && c986_inl1_inl49);
  assign c2901 = (c2895 && c848_inl51);
  assign c2902 = (c2900 && c988_inl1_inl49);
  assign c2903 = (c2900 && !c988_inl1_inl49);
  assign c2904 = (c2876 && !c986_inl1_inl49);
  assign c2905 = (c2901 && !c994_inl1_inl1_inl51);
  assign c2906 = ((c2904 || c2902) && c986_inl2_inl49);
  assign c2907 = (c2901 && !c985_inl2_inl1_inl51);
  assign c2908 = (c2906 && c988_inl2_inl49);
  assign c2909 = (c2906 && !c988_inl2_inl49);
  assign c2910 = ((c2904 || c2902) && !c986_inl2_inl49);
  assign c2911 = (c2901 && !c985_inl3_inl1_inl51);
  assign c2912 = (c2901 && c851_inl51);
  assign c2913 = ((c2910 || c2908) && c973_inl49);
  assign c2914 = (c2895 && !c848_inl51);
  assign c2915 = (c2901 && !c851_inl51);
  assign c2916 = (((c2914 || c2915) || c2912) && c853_inl51);
  assign c2917 = (c2916 && c856_inl51);
  assign c2918 = (c2916 && !c856_inl51);
  assign c2919 = (c2917 && c857_inl51);
  assign c2920 = (c2917 && !c857_inl51);
  assign c2921 = (c2919 && !c994_inl1_inl5_inl51);
  assign c2922 = (c2920 && !c994_inl1_inl8_inl51);
  assign c2923 = (c2919 && !c985_inl2_inl5_inl51);
  assign c2924 = (c2920 && !c985_inl2_inl8_inl51);
  assign c2925 = (c2919 && !c985_inl3_inl5_inl51);
  assign c2926 = (c2920 && !c985_inl3_inl8_inl51);
  assign c2927 = (c2919 && !c994_inl1_inl6_inl51);
  assign c2928 = (c2919 && !c985_inl2_inl6_inl51);
  assign c2929 = (c2919 && !c985_inl3_inl6_inl51);
  assign c2930 = (c2919 && !c994_inl1_inl7_inl51);
  assign c2931 = (c2919 && !c985_inl2_inl7_inl51);
  assign c2932 = (c2920 && c985_inl3_inl8_inl51);
  assign c2933 = (c2919 && c985_inl3_inl7_inl51);
  assign c2934 = (c2919 && !c985_inl3_inl7_inl51);
  assign c2935 = (((c2918 || c2932) || c2933) && !c994_inl1_inl9_inl51);
  assign c2936 = (((c2918 || c2932) || c2933) && !c985_inl2_inl9_inl51);
  assign c2937 = (((c2918 || c2932) || c2933) && !c985_inl3_inl9_inl51);
  assign c2938 = (((c2914 || c2915) || c2912) && !c853_inl51);
  assign c2939 = ((c2918 || c2932) || c2933);
  assign c2940 = ((c2938 || c2939) && c860_inl51);
  assign c2941 = ((c2938 || c2939) && !c860_inl51);
  assign c2942 = ((c2941 || c2940) && c862_inl51);
  assign c2943 = ((c2941 || c2940) && !c862_inl51);
  assign c2944 = ((c2943 || c2942) && c864_inl51);
  assign c2945 = ((c2943 || c2942) && c1084_inl51);
  assign c2946 = ((c2943 || c2942) && c1085_inl51);
  assign c2947 = ((c2943 || c2942) && c1086_inl51);
  assign c2948 = ((c2943 || c2942) && c1087_inl51);
  assign c2949 = ((c2943 || c2942) && c1088_inl51);
  assign c2950 = ((c2943 || c2942) && c1089_inl51);
  assign c2951 = ((c2943 || c2942) && c1090_inl51);
  assign c2952 = ((((((((c2951 || c2946) || c2944) || c2945) || c2950) || c2949) || c2948) || c2947) && c878_inl51);
  assign c2953 = ((((((((c2951 || c2946) || c2944) || c2945) || c2950) || c2949) || c2948) || c2947) && !c878_inl51);
  assign c2954 = ((c2953 || c2952) && c880_inl51);
  assign c2955 = ((c2953 || c2952) && c1091_inl51);
  assign c2956 = ((c2953 || c2952) && c1092_inl51);
  assign c2957 = ((c2953 || c2952) && c1093_inl51);
  assign c2958 = ((c2953 || c2952) && c1094_inl51);
  assign c2959 = ((c2953 || c2952) && c1095_inl51);
  assign c2960 = ((c2953 || c2952) && c1096_inl51);
  assign c2961 = ((c2953 || c2952) && c1097_inl51);
  assign c2962 = ((c2953 || c2952) && c1098_inl51);
  assign c2963 = ((c2953 || c2952) && c1099_inl51);
  assign c2964 = ((c2953 || c2952) && c1100_inl51);
  assign c2965 = ((c2953 || c2952) && c1101_inl51);
  assign c2966 = ((c2953 || c2952) && c1102_inl51);
  assign c2967 = ((c2953 || c2952) && c1103_inl51);
  assign c2968 = ((c2953 || c2952) && c1104_inl51);
  assign c2969 = ((c2953 || c2952) && c1105_inl51);
  assign c2970 = ((((((((((((((((c2969 || c2959) || c2954) || c2967) || c2958) || c2957) || c2960) || c2961) || c2966) || c2963) || c2965) || c2968) || c2964) || c2956) || c2962) || c2955) && c910_inl51);
  assign c2971 = ((((((((((((((((c2969 || c2959) || c2954) || c2967) || c2958) || c2957) || c2960) || c2961) || c2966) || c2963) || c2965) || c2968) || c2964) || c2956) || c2962) || c2955) && !c910_inl51);
  assign c848_inl51 = (t847_inl51 == 1);
  assign c851_inl51 = (t850_inl51 == 13);
  assign c853_inl51 = (t852_inl51 == 1);
  assign c854_inl51 = (stack0_top2 > 0);
  assign c855_inl51 = (stack0_top2 < 128);
  assign c856_inl51 = (c854_inl51 && c855_inl51);
  assign c857_inl51 = (stack0_top2 == 8);
  assign c860_inl51 = (t859_inl51 == 1);
  assign c862_inl51 = (t861_inl51 == 2);
  assign c864_inl51 = (t863_inl51 == -1);
  assign c866_inl51 = (t865_inl51 == -2);
  assign c868_inl51 = (t867_inl51 == -3);
  assign c870_inl51 = (t869_inl51 == -4);
  assign c872_inl51 = (t871_inl51 == -5);
  assign c874_inl51 = (t873_inl51 == -6);
  assign c876_inl51 = (t875_inl51 == -7);
  assign c878_inl51 = (t877_inl51 == -8);
  assign c880_inl51 = (t879_inl51 == -1);
  assign c882_inl51 = (t881_inl51 == -2);
  assign c884_inl51 = (t883_inl51 == -3);
  assign c886_inl51 = (t885_inl51 == -4);
  assign c888_inl51 = (t887_inl51 == -5);
  assign c890_inl51 = (t889_inl51 == -6);
  assign c892_inl51 = (t891_inl51 == -7);
  assign c894_inl51 = (t893_inl51 == -8);
  assign c896_inl51 = (t895_inl51 == -9);
  assign c898_inl51 = (t897_inl51 == -10);
  assign c900_inl51 = (t899_inl51 == -11);
  assign c902_inl51 = (t901_inl51 == -12);
  assign c904_inl51 = (t903_inl51 == -13);
  assign c906_inl51 = (t905_inl51 == -14);
  assign c908_inl51 = (t907_inl51 == -15);
  assign c910_inl51 = (t909_inl51 == 1);
  assign c914 = (ip2 < 16384);
  assign c915 = (opcode3 <= 30);
  assign c916 = (opcode3 == 0);
  assign c917 = (opcode3 == 1);
  assign c918 = (opcode3 == 2);
  assign c919 = (opcode3 == 3);
  assign c920 = (opcode3 == 4);
  assign c921 = (opcode3 == 5);
  assign c922 = (opcode3 == 6);
  assign c923 = (opcode3 == 7);
  assign c924 = (opcode3 == 8);
  assign c925 = (opcode3 == 9);
  assign c926 = (opcode3 == 10);
  assign c927 = (opcode3 == 11);
  assign c928 = (opcode3 == 12);
  assign c929 = (opcode3 == 13);
  assign c930 = (opcode3 == 14);
  assign c931 = (opcode3 == 15);
  assign c932 = (opcode3 == 16);
  assign c933 = (opcode3 == 17);
  assign c934 = (opcode3 == 18);
  assign c935 = (opcode3 == 19);
  assign c936 = (opcode3 == 20);
  assign c937 = (opcode3 == 21);
  assign c938 = (opcode3 == 22);
  assign c939 = (opcode3 == 23);
  assign c940 = (opcode3 == 24);
  assign c941 = (opcode3 == 25);
  assign c942 = (opcode3 == 26);
  assign c943 = (opcode3 == 27);
  assign c944 = (opcode3 == 28);
  assign c945 = (opcode3 == 29);
  assign c946 = (opcode3 == 30);
  assign c950 = (stack0_top9 != 0);
  assign c951 = (stack0_top9 > -1);
  assign c952 = (c950 && c951);
  assign c955 = (stack0_second2 > stack0_top2);
  assign c957 = (stack0_second2 < stack0_top2);
  assign c959 = (stack0_second2 != stack0_top2);
  assign c961 = (stack0_second2 == stack0_top2);
  assign c964 = (stack0_top2 == 0);
  assign c967 = (t966 == 0);
  assign c973_inl49 = (i_inl493 < t486_inl49);
  assign c974_inl49 = (abs_a_inl493 >= abs_b_inl494);
  assign c975_inl49 = (t970_inl49 != 0);
  assign c977_inl49 = (t976_inl49 != 0);
  assign c985_inl2_inl1_inl51 = (cmd_reply_inl2_inl1_inl51 == 2147483650);
  assign c985_inl2_inl5_inl51 = (cmd_reply_inl2_inl5_inl51 == 2147483649);
  assign c985_inl2_inl6_inl51 = (cmd_reply_inl2_inl6_inl51 == 2147483649);
  assign c985_inl2_inl7_inl51 = (cmd_reply_inl2_inl7_inl51 == 2147483649);
  assign c985_inl2_inl8_inl51 = (cmd_reply_inl2_inl8_inl51 == 2147483649);
  assign c985_inl2_inl9_inl51 = (cmd_reply_inl2_inl9_inl51 == 2147483651);
  assign c985_inl3_inl1_inl51 = (cmd_reply_inl3_inl1_inl51 == 2147483648);
  assign c985_inl3_inl5_inl51 = (cmd_reply_inl3_inl5_inl51 == 2147483648);
  assign c985_inl3_inl6_inl51 = (cmd_reply_inl3_inl6_inl51 == 2147483648);
  assign c985_inl3_inl7_inl51 = (cmd_reply_inl3_inl7_inl51 == 2147483648);
  assign c985_inl3_inl8_inl51 = (cmd_reply_inl3_inl8_inl51 == 2147483648);
  assign c985_inl3_inl9_inl51 = (cmd_reply_inl3_inl9_inl51 == 2147483648);
  assign c986_inl1_inl49 = (i_inl1_inl493 < 31);
  assign c986_inl2_inl49 = (i_inl2_inl493 < 31);
  assign c988_inl1_inl49 = (t987_inl1_inl49 != 0);
  assign c988_inl2_inl49 = (t987_inl2_inl49 != 0);
  assign c994_inl1_inl1_inl51 = (t993_inl1_inl1_inl51 == 0);
  assign c994_inl1_inl5_inl51 = (t993_inl1_inl5_inl51 == 0);
  assign c994_inl1_inl6_inl51 = (t993_inl1_inl6_inl51 == 0);
  assign c994_inl1_inl7_inl51 = (t993_inl1_inl7_inl51 == 0);
  assign c994_inl1_inl8_inl51 = (t993_inl1_inl8_inl51 == 0);
  assign c994_inl1_inl9_inl51 = (t993_inl1_inl9_inl51 == 0);
  assign c_bit_inl494 = (c_bit_inl493 | 2147483648);
  assign c_bit_inl495 = c2299 ? c_bit_inl494 : ((c2296 || c2294) && !c977_inl49) ? c_bit_inl493 : 'bz;
  assign c_bit_inl496 = (c_bit_inl493 << 1);
  assign c_bit_inl497 = (c_bit_inl496 | 1);
  assign c_bit_inl498 = (c_bit_inl493 << 1);
  assign c_bit_inl499 = c2292 ? c_bit_inl497 : c2293 ? c_bit_inl498 : 'bz;
  assign cmd_reply_inl1_inl1_inl51 = (t992_inl1_inl1_inl51 & 4294967295);
  assign cmd_reply_inl1_inl5_inl51 = (t992_inl1_inl5_inl51 & 4294967295);
  assign cmd_reply_inl1_inl6_inl51 = (t992_inl1_inl6_inl51 & 4294967295);
  assign cmd_reply_inl1_inl7_inl51 = (t992_inl1_inl7_inl51 & 4294967295);
  assign cmd_reply_inl1_inl8_inl51 = (t992_inl1_inl8_inl51 & 4294967295);
  assign cmd_reply_inl1_inl9_inl51 = (t992_inl1_inl9_inl51 & 4294967295);
  assign cmd_reply_inl2_inl1_inl51 = (t983_inl2_inl1_inl51 & 4294967295);
  assign cmd_reply_inl2_inl5_inl51 = (t983_inl2_inl5_inl51 & 4294967295);
  assign cmd_reply_inl2_inl6_inl51 = (t983_inl2_inl6_inl51 & 4294967295);
  assign cmd_reply_inl2_inl7_inl51 = (t983_inl2_inl7_inl51 & 4294967295);
  assign cmd_reply_inl2_inl8_inl51 = (t983_inl2_inl8_inl51 & 4294967295);
  assign cmd_reply_inl2_inl9_inl51 = (t983_inl2_inl9_inl51 & 4294967295);
  assign cmd_reply_inl3_inl1_inl51 = (t983_inl3_inl1_inl51 & 4294967295);
  assign cmd_reply_inl3_inl5_inl51 = (t983_inl3_inl5_inl51 & 4294967295);
  assign cmd_reply_inl3_inl6_inl51 = (t983_inl3_inl6_inl51 & 4294967295);
  assign cmd_reply_inl3_inl7_inl51 = (t983_inl3_inl7_inl51 & 4294967295);
  assign cmd_reply_inl3_inl8_inl51 = (t983_inl3_inl8_inl51 & 4294967295);
  assign cmd_reply_inl3_inl9_inl51 = (t983_inl3_inl9_inl51 & 4294967295);
  assign find_zero_len_result2_inl494 = c2284 ? n_inl2_inl493 : (c2177 || c2256) ? 0 : 'bz;
  assign i_inl1_inl494 = (i_inl1_inl493 + 1);
  assign i_inl2_inl494 = (i_inl2_inl493 + 1);
  assign i_inl494 = (i_inl493 + 1);
  assign ip10 = (ip2 + 1);
  assign ip11 = (t956 - 1);
  assign ip12 = (ip2 + 1);
  assign ip13 = (t958 - 1);
  assign ip14 = (ip2 + 1);
  assign ip15 = (t960 - 1);
  assign ip16 = (ip2 + 1);
  assign ip17 = (t962 - 1);
  assign ip20 = (t968 - 1);
  assign ip21 = (c2157 && c916) ? ip2 : c2159 ? ip3 : c2160 ? ip2 : c2161 ? ip2 : c2162 ? ip2 : c2163 ? ip2 : c2164 ? ip2 : c2246 ? ip5 : c2247 ? ip6 : c2166 ? ip8 : c2167 ? address0_top2 : c2168 ? t2660 : c2169 ? t2670 : c2170 ? t2680 : c2171 ? t2690 : c2172 ? ip2 : c2173 ? ip2 : c2174 ? ip2 : c2175 ? ip2 : c2176 ? ip2 : (c2286 || c2284) ? ip2 : c2178 ? ip2 : c2179 ? ip2 : c2180 ? ip2 : c2181 ? ip2 : c2182 ? ip2 : c2212 ? address0_top2 : (c2183 && !c964) ? ip2 : c2184 ? ip2 : c2185 ? ip2 : c2186 ? ip2 : c2187 ? ip2 : (c2361 || c2360) ? ip_inl514 : (c2188 && !c967) ? ip2 : (c2157 && c1136) ? ip2 : c2158 ? ip20 : 'bz;
  assign ip22 = (ip21 + 1);
  assign ip3 = (ip2 + 1);
  assign ip4 = (ip2 + 1);
  assign ip5 = (t953 - 1);
  assign ip6 = (ip2 + 1);
  assign ip7 = (ip2 + 1);
  assign ip8 = (t954 - 1);
  assign ip_inl514 = c2344 ? ip2 : c2345 ? ip2 : c2346 ? ip2 : c2347 ? ip2 : c2348 ? ip2 : c2349 ? ip2 : c2350 ? ip2 : c2351 ? ip2 : c2352 ? 16384 : c2353 ? ip2 : c2354 ? ip2 : c2355 ? ip2 : c2356 ? ip2 : c2357 ? ip2 : c2358 ? ip2 : ((c2343 || c2342) && c1105_inl51) ? ip2 : 'bz;
  assign n_inl1_inl494 = (n_inl1_inl493 + 1);
  assign n_inl2_inl494 = (n_inl2_inl493 + 1);
  assign retro_divmod_result492[0] = array995_inl49[0];
  assign retro_divmod_result492[1] = array995_inl49[1];
  assign stack0_pos10 = (stack0_pos9 - 1);
  assign stack0_pos11 = (stack0_pos2 - 1);
  assign stack0_pos12 = (stack0_pos11 - 1);
  assign stack0_pos13 = (stack0_pos2 - 1);
  assign stack0_pos14 = (stack0_pos13 - 1);
  assign stack0_pos15 = (stack0_pos2 - 1);
  assign stack0_pos16 = (stack0_pos15 - 1);
  assign stack0_pos17 = (stack0_pos2 - 1);
  assign stack0_pos18 = (stack0_pos17 - 1);
  assign stack0_pos19 = (stack0_pos2 - 1);
  assign stack0_pos20 = (stack0_pos2 - 1);
  assign stack0_pos21 = (stack0_pos2 - 1);
  assign stack0_pos22 = (stack0_pos2 - 1);
  assign stack0_pos23 = (stack0_pos2 - 1);
  assign stack0_pos24 = (stack0_pos2 - 1);
  assign stack0_pos25 = (stack0_pos2 - 1);
  assign stack0_pos26 = (stack0_pos2 - 1);
  assign stack0_pos27 = (stack0_pos2 - 1);
  assign stack0_pos28 = (stack0_pos2 - 1);
  assign stack0_pos29 = (stack0_pos28 - 1);
  assign stack0_pos30 = (stack0_pos2 - 1);
  assign stack0_pos31 = (stack0_pos2 - 1);
  assign stack0_pos32 = (stack0_pos2 - 1);
  assign stack0_pos33 = (c2300 && c985_inl3_inl7_inl51) ? stack0_pos30 : (c2301 && c985_inl3_inl8_inl51) ? stack0_pos31 : c2298 ? stack0_pos32 : 'bz;
  assign stack0_pos34 = ((c2298 || c2322) || c2323) ? stack0_pos33 : (((c2290 || c2291) || c2288) && !c853_inl51) ? stack0_pos2 : 'bz;
  assign stack0_pos35 = (c2157 && c916) ? stack0_pos2 : c2159 ? stack0_pos3 : c2160 ? stack0_pos4 : c2161 ? stack0_pos5 : c2162 ? stack0_pos2 : c2163 ? stack0_pos6 : c2164 ? stack0_pos7 : c2246 ? stack0_pos2 : c2247 ? stack0_pos8 : c2166 ? stack0_pos2 : c2167 ? stack0_pos2 : c2168 ? stack0_pos10 : c2169 ? stack0_pos12 : c2170 ? stack0_pos14 : c2171 ? stack0_pos16 : c2172 ? stack0_pos2 : c2173 ? stack0_pos18 : c2174 ? stack0_pos19 : c2175 ? stack0_pos20 : c2176 ? stack0_pos21 : (c2286 || c2284) ? stack0_pos2 : c2178 ? stack0_pos22 : c2179 ? stack0_pos23 : c2180 ? stack0_pos24 : c2181 ? stack0_pos25 : c2182 ? stack0_pos26 : c2212 ? stack0_pos27 : (c2183 && !c964) ? stack0_pos2 : c2184 ? stack0_pos2 : c2185 ? stack0_pos2 : c2186 ? stack0_pos2 : c2187 ? stack0_pos29 : (c2361 || c2360) ? stack0_pos34 : (c2188 && !c967) ? stack0_pos2 : (c2157 && c1136) ? stack0_pos2 : c2158 ? stack0_pos2 : 'bz;
  assign stack0_pos3 = (stack0_pos2 + 1);
  assign stack0_pos4 = (stack0_pos2 + 1);
  assign stack0_pos5 = (stack0_pos2 - 1);
  assign stack0_pos6 = (stack0_pos2 - 1);
  assign stack0_pos7 = (stack0_pos2 + 1);
  assign stack0_pos8 = (stack0_pos2 - 1);
  assign stack0_pos9 = (stack0_pos2 - 1);
  assign stack0_second23 = retro_divmod_result492[1];
  assign stack0_second35 = (c2300 && c985_inl3_inl7_inl51) ? stack0_second32 : (c2301 && c985_inl3_inl8_inl51) ? stack0_second33 : c2298 ? stack0_second34 : 'bz;
  assign stack0_second36 = ((c2298 || c2322) || c2323) ? stack0_second35 : (((c2290 || c2291) || c2288) && !c853_inl51) ? stack0_second2 : 'bz;
  assign stack0_second37 = (c2157 && c916) ? stack0_second2 : c2159 ? stack0_top2 : c2160 ? stack0_top2 : c2161 ? stack0_second5 : c2162 ? stack0_top2 : c2163 ? stack0_second7 : c2164 ? stack0_top2 : c2246 ? stack0_second2 : c2247 ? stack0_second9 : c2166 ? stack0_second2 : c2167 ? stack0_second2 : c2168 ? stack0_second11 : c2169 ? stack0_second13 : c2170 ? stack0_second15 : c2171 ? stack0_second17 : c2172 ? stack0_second2 : c2173 ? stack0_second19 : c2174 ? stack0_second20 : c2175 ? stack0_second21 : c2176 ? stack0_second22 : (c2286 || c2284) ? stack0_second23 : c2178 ? stack0_second24 : c2179 ? stack0_second25 : c2180 ? stack0_second26 : c2181 ? stack0_second27 : c2182 ? stack0_second28 : c2212 ? stack0_second29 : (c2183 && !c964) ? stack0_second2 : c2184 ? stack0_second2 : c2185 ? stack0_second2 : c2186 ? stack0_second2 : c2187 ? stack0_second31 : (c2361 || c2360) ? stack0_second36 : (c2188 && !c967) ? stack0_second2 : (c2157 && c1136) ? stack0_second2 : c2158 ? stack0_second2 : 'bz;
  assign stack0_top23 = (stack0_second2 + stack0_top2);
  assign stack0_top25 = (stack0_second2 - stack0_top2);
  assign stack0_top27 = (stack0_second2 * stack0_top2);
  assign stack0_top28 = retro_divmod_result492[0];
  assign stack0_top30 = (stack0_second2 & stack0_top2);
  assign stack0_top32 = (stack0_second2 | stack0_top2);
  assign stack0_top34 = (stack0_second2 ^ stack0_top2);
  assign stack0_top36 = (stack0_second2 << stack0_top2);
  assign stack0_top38 = (stack0_second2 >>> stack0_top2);
  assign stack0_top40 = (stack0_top2 + 1);
  assign stack0_top41 = (stack0_top2 - 1);
  assign stack0_top49 = ((c2298 || c2322) || c2323) ? stack0_second2 : (((c2290 || c2291) || c2288) && !c853_inl51) ? stack0_top2 : 'bz;
  assign stack0_top50 = (c2157 && c916) ? stack0_top2 : c2159 ? t947 : c2160 ? stack0_top2 : c2161 ? stack0_second2 : c2162 ? stack0_second2 : c2163 ? stack0_second2 : c2164 ? address0_top2 : c2246 ? stack0_top9 : c2247 ? stack0_second2 : c2166 ? stack0_top2 : c2167 ? stack0_top2 : c2168 ? stack0_second10 : c2169 ? stack0_second12 : c2170 ? stack0_second14 : c2171 ? stack0_second16 : c2172 ? stack0_top19 : c2173 ? stack0_second18 : c2174 ? stack0_top23 : c2175 ? stack0_top25 : c2176 ? stack0_top27 : (c2286 || c2284) ? stack0_top28 : c2178 ? stack0_top30 : c2179 ? stack0_top32 : c2180 ? stack0_top34 : c2181 ? stack0_top36 : c2182 ? stack0_top38 : c2212 ? stack0_second2 : (c2183 && !c964) ? stack0_top2 : c2184 ? stack0_top40 : c2185 ? stack0_top41 : c2186 ? stack0_top42 : c2187 ? stack0_second30 : (c2361 || c2360) ? stack0_top49 : (c2188 && !c967) ? stack0_top2 : (c2157 && c1136) ? stack0_top2 : c2158 ? stack0_top2 : 'bz;
  assign stack0_top9 = (stack0_top2 - 1);
  assign t2660 = c2277 ? ip11 : (c2168 && !c955) ? ip10 : 'bz;
  assign t2670 = c2278 ? ip13 : (c2169 && !c957) ? ip12 : 'bz;
  assign t2680 = c2279 ? ip15 : (c2170 && !c959) ? ip14 : 'bz;
  assign t2690 = c2280 ? ip17 : (c2171 && !c961) ? ip16 : 'bz;
  assign t486_inl49 = (find_zero_len_result2_inl494 + 1);
  assign t843_inl3 = (stack0_pos2 - 2);
  assign t843_inl4 = (stack0_pos2 - 2);
  assign t843_inl5 = (address0_pos2 - 2);
  assign t843_inl6 = (stack0_pos2 - 2);
  assign t843_inl7 = (address0_pos2 - 2);
  assign t846_inl10 = (address0_pos4 - 2);
  assign t846_inl11 = (stack0_pos8 - 2);
  assign t846_inl12 = (address0_pos5 - 2);
  assign t846_inl13 = (stack0_pos9 - 2);
  assign t846_inl14 = (stack0_pos10 - 2);
  assign t846_inl15 = (stack0_pos11 - 2);
  assign t846_inl16 = (stack0_pos12 - 2);
  assign t846_inl17 = (stack0_pos13 - 2);
  assign t846_inl18 = (stack0_pos14 - 2);
  assign t846_inl19 = (stack0_pos15 - 2);
  assign t846_inl20 = (stack0_pos16 - 2);
  assign t846_inl21 = (stack0_pos17 - 2);
  assign t846_inl22 = (stack0_pos18 - 2);
  assign t846_inl23 = (stack0_pos19 - 2);
  assign t846_inl24 = (stack0_pos20 - 2);
  assign t846_inl25 = (stack0_pos21 - 2);
  assign t846_inl26 = (stack0_pos22 - 2);
  assign t846_inl27 = (stack0_pos23 - 2);
  assign t846_inl28 = (stack0_pos24 - 2);
  assign t846_inl29 = (stack0_pos25 - 2);
  assign t846_inl2_inl51 = (stack0_pos30 - 2);
  assign t846_inl30 = (stack0_pos26 - 2);
  assign t846_inl31 = (stack0_pos27 - 2);
  assign t846_inl32 = (address0_pos6 - 2);
  assign t846_inl33 = (stack0_pos28 - 2);
  assign t846_inl34 = (stack0_pos29 - 2);
  assign t846_inl3_inl51 = (stack0_pos31 - 2);
  assign t846_inl4_inl51 = (stack0_pos32 - 2);
  assign t846_inl8 = (stack0_pos5 - 2);
  assign t846_inl9 = (stack0_pos6 - 2);
  assign t969_inl49 = (stack0_second2 & 2147483648);
  assign t970_inl49 = t969_inl49 ? 1 : 0;
  assign t971_inl49 = (stack0_top2 & 2147483648);
  assign t972_inl49 = t971_inl49 ? 1 : 0;
  assign t976_inl49 = (t970_inl49 ^ t972_inl49);
  assign t987_inl1_inl49 = (test_bit_inl1_inl493 & x_inl1_inl49);
  assign t987_inl2_inl49 = (test_bit_inl2_inl493 & x_inl2_inl49);
  assign t993_inl1_inl1_inl51 = (cmd_reply_inl1_inl1_inl51 & 2147483648);
  assign t993_inl1_inl5_inl51 = (cmd_reply_inl1_inl5_inl51 & 2147483648);
  assign t993_inl1_inl6_inl51 = (cmd_reply_inl1_inl6_inl51 & 2147483648);
  assign t993_inl1_inl7_inl51 = (cmd_reply_inl1_inl7_inl51 & 2147483648);
  assign t993_inl1_inl8_inl51 = (cmd_reply_inl1_inl8_inl51 & 2147483648);
  assign t993_inl1_inl9_inl51 = (cmd_reply_inl1_inl9_inl51 & 2147483648);
  assign test_bit_inl1_inl494 = (test_bit_inl1_inl493 >>> 1);
  assign test_bit_inl2_inl494 = (test_bit_inl2_inl493 >>> 1);
  assign x_inl1_inl49 = abs_a_inl492;
  assign x_inl2_inl49 = abs_b_inl492;
  //combinations: array996
  assign _stack_len = array996_ram_len;
  assign _stack_q = array996_ram_q;
  assign array996_ram_addr = _stack_addr;
  assign array996_ram_d = _stack_d;
  assign array996_ram_we = _stack_we;
  //combinations: array997
  assign _address_len = array997_ram_len;
  assign _address_q = array997_ram_q;
  assign array997_ram_addr = _address_addr;
  assign array997_ram_d = _address_d;
  assign array997_ram_we = _address_we;
  //combinations: in_io_ports
  assign io_ports_len = retro_main_in_io_ports_len;
  assign io_ports_q = retro_main_in_io_ports_q;
  assign retro_main_in_io_ports_addr = io_ports_addr;
  assign retro_main_in_io_ports_d = io_ports_d;
  assign retro_main_in_io_ports_req = io_ports_req;
  assign retro_main_in_io_ports_we = io_ports_we;
  //combinations: in_memory
  assign memory_len = retro_main_in_memory_len;
  assign memory_q = retro_main_in_memory_q;
  assign retro_main_in_memory_addr = memory_addr;
  assign retro_main_in_memory_d = memory_d;
  assign retro_main_in_memory_req = memory_req;
  assign retro_main_in_memory_we = memory_we;
  //sub modules
  //array996 instance
  BidirectionalSinglePortRam#(
    .DATA_WIDTH(32),
    .ADDR_WIDTH(8),
    .RAM_LENGTH(128)
    )
    array996(
      .clk(clk),
      .rst(rst),
      .ram_addr(array996_ram_addr),
      .ram_d(array996_ram_d),
      .ram_we(array996_ram_we),
      .ram_q(array996_ram_q),
      .ram_len(array996_ram_len)
    );
  //array997 instance
  BidirectionalSinglePortRam#(
    .DATA_WIDTH(32),
    .ADDR_WIDTH(11),
    .RAM_LENGTH(1024)
    )
    array997(
      .clk(clk),
      .rst(rst),
      .ram_addr(array997_ram_addr),
      .ram_d(array997_ram_d),
      .ram_we(array997_ram_we),
      .ram_q(array997_ram_q),
      .ram_len(array997_ram_len)
    );
  
  
  always @(posedge clk) begin
    if (rst) begin
      _address_addr <= 0;
      _address_d <= 0;
      _address_req <= 0;
      _address_we <= 0;
      _stack_addr <= 0;
      _stack_d <= 0;
      _stack_req <= 0;
      _stack_we <= 0;
      a6 <= 0;
      abs_a_inl493 <= 0;
      abs_b_inl494 <= 0;
      address0_pos2 <= 0;
      address0_second2 <= 0;
      address0_second4 <= 0;
      address0_second5 <= 0;
      address0_second6 <= 0;
      address0_top2 <= 0;
      b6 <= 0;
      c_bit_inl493 <= 0;
      char_c_inl1_inl51 <= 0;
      i_inl1_inl493 <= 0;
      i_inl2_inl493 <= 0;
      i_inl493 <= 0;
      io_ports_addr <= 0;
      io_ports_d <= 0;
      io_ports_req <= 0;
      io_ports_we <= 0;
      ip2 <= 0;
      memory_addr <= 0;
      memory_d <= 0;
      memory_req <= 0;
      memory_we <= 0;
      n_inl1_inl493 <= 0;
      n_inl2_inl493 <= 0;
      opcode3 <= 0;
      stack0_pos2 <= 0;
      stack0_second10 <= 0;
      stack0_second11 <= 0;
      stack0_second12 <= 0;
      stack0_second13 <= 0;
      stack0_second14 <= 0;
      stack0_second15 <= 0;
      stack0_second16 <= 0;
      stack0_second17 <= 0;
      stack0_second18 <= 0;
      stack0_second19 <= 0;
      stack0_second20 <= 0;
      stack0_second21 <= 0;
      stack0_second22 <= 0;
      stack0_second24 <= 0;
      stack0_second25 <= 0;
      stack0_second26 <= 0;
      stack0_second27 <= 0;
      stack0_second28 <= 0;
      stack0_second29 <= 0;
      stack0_second2 <= 0;
      stack0_second30 <= 0;
      stack0_second31 <= 0;
      stack0_second32 <= 0;
      stack0_second33 <= 0;
      stack0_second34 <= 0;
      stack0_second5 <= 0;
      stack0_second7 <= 0;
      stack0_second9 <= 0;
      stack0_top19 <= 0;
      stack0_top2 <= 0;
      stack0_top42 <= 0;
      t11 <= 0;
      t847_inl51 <= 0;
      t850_inl51 <= 0;
      t852_inl51 <= 0;
      t859_inl51 <= 0;
      t861_inl51 <= 0;
      t863_inl51 <= 0;
      t865_inl51 <= 0;
      t867_inl51 <= 0;
      t869_inl51 <= 0;
      t871_inl51 <= 0;
      t873_inl51 <= 0;
      t875_inl51 <= 0;
      t877_inl51 <= 0;
      t879_inl51 <= 0;
      t881_inl51 <= 0;
      t883_inl51 <= 0;
      t885_inl51 <= 0;
      t887_inl51 <= 0;
      t889_inl51 <= 0;
      t891_inl51 <= 0;
      t893_inl51 <= 0;
      t895_inl51 <= 0;
      t897_inl51 <= 0;
      t899_inl51 <= 0;
      t901_inl51 <= 0;
      t903_inl51 <= 0;
      t905_inl51 <= 0;
      t907_inl51 <= 0;
      t909_inl51 <= 0;
      t947 <= 0;
      t953 <= 0;
      t954 <= 0;
      t956 <= 0;
      t958 <= 0;
      t960 <= 0;
      t962 <= 0;
      t966 <= 0;
      t968 <= 0;
      t983_inl2_inl1_inl51 <= 0;
      t983_inl2_inl5_inl51 <= 0;
      t983_inl2_inl6_inl51 <= 0;
      t983_inl2_inl7_inl51 <= 0;
      t983_inl2_inl8_inl51 <= 0;
      t983_inl2_inl9_inl51 <= 0;
      t983_inl3_inl1_inl51 <= 0;
      t983_inl3_inl5_inl51 <= 0;
      t983_inl3_inl6_inl51 <= 0;
      t983_inl3_inl7_inl51 <= 0;
      t983_inl3_inl8_inl51 <= 0;
      t983_inl3_inl9_inl51 <= 0;
      t992_inl1_inl1_inl51 <= 0;
      t992_inl1_inl5_inl51 <= 0;
      t992_inl1_inl6_inl51 <= 0;
      t992_inl1_inl7_inl51 <= 0;
      t992_inl1_inl8_inl51 <= 0;
      t992_inl1_inl9_inl51 <= 0;
      test_bit_inl1_inl493 <= 0;
      test_bit_inl2_inl493 <= 0;
      retro_main_state <= retro_main_b1_INIT;
    end else begin //if (rst)
      case(retro_main_state)
      retro_main_b1_INIT: begin
        retro_main_valid <= 0;
        if (retro_main_ready == 1) begin
          _address_addr <= 0;
          _address_we <= 1;
          _address_req <= 1;
          _address_d <= 0;
          _stack_addr <= 0;
          _stack_we <= 1;
          _stack_req <= 1;
          _stack_d <= 0;
          array998[0] <= 0;
          array998[1] <= 0;
          array998[2] <= 0;
          array998[3] <= 0;
          array998[4] <= 0;
          array998[5] <= 0;
          array998[6] <= 0;
          array998[7] <= 0;
          array998[8] <= 0;
          array998[9] <= 0;
          array998[10] <= 0;
          array998[11] <= 0;
          address0_pos2 <= 0;
          address0_second2 <= 0;
          address0_top2 <= 0;
          ip2 <= 0;
          stack0_pos2 <= 0;
          stack0_second2 <= 0;
          stack0_top2 <= 0;
          retro_main_state <= retro_main_b1_S1;
        end
      end
      retro_main_b1_S1: begin
        _address_addr <= 1;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 1;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S2;
      end
      retro_main_b1_S2: begin
        _address_addr <= 2;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 2;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S3;
      end
      retro_main_b1_S3: begin
        _address_addr <= 3;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 3;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S4;
      end
      retro_main_b1_S4: begin
        _address_addr <= 4;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 4;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S5;
      end
      retro_main_b1_S5: begin
        _address_addr <= 5;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 5;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S6;
      end
      retro_main_b1_S6: begin
        _address_addr <= 6;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 6;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S7;
      end
      retro_main_b1_S7: begin
        _address_addr <= 7;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 7;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S8;
      end
      retro_main_b1_S8: begin
        _address_addr <= 8;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 8;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S9;
      end
      retro_main_b1_S9: begin
        _address_addr <= 9;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 9;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S10;
      end
      retro_main_b1_S10: begin
        _address_addr <= 10;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 10;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S11;
      end
      retro_main_b1_S11: begin
        _address_addr <= 11;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 11;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S12;
      end
      retro_main_b1_S12: begin
        _address_addr <= 12;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 12;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S13;
      end
      retro_main_b1_S13: begin
        _address_addr <= 13;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 13;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S14;
      end
      retro_main_b1_S14: begin
        _address_addr <= 14;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 14;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S15;
      end
      retro_main_b1_S15: begin
        _address_addr <= 15;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 15;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S16;
      end
      retro_main_b1_S16: begin
        _address_addr <= 16;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 16;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S17;
      end
      retro_main_b1_S17: begin
        _address_addr <= 17;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 17;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S18;
      end
      retro_main_b1_S18: begin
        _address_addr <= 18;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 18;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S19;
      end
      retro_main_b1_S19: begin
        _address_addr <= 19;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 19;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S20;
      end
      retro_main_b1_S20: begin
        _address_addr <= 20;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 20;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S21;
      end
      retro_main_b1_S21: begin
        _address_addr <= 21;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 21;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S22;
      end
      retro_main_b1_S22: begin
        _address_addr <= 22;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 22;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S23;
      end
      retro_main_b1_S23: begin
        _address_addr <= 23;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 23;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S24;
      end
      retro_main_b1_S24: begin
        _address_addr <= 24;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 24;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S25;
      end
      retro_main_b1_S25: begin
        _address_addr <= 25;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 25;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S26;
      end
      retro_main_b1_S26: begin
        _address_addr <= 26;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 26;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S27;
      end
      retro_main_b1_S27: begin
        _address_addr <= 27;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 27;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S28;
      end
      retro_main_b1_S28: begin
        _address_addr <= 28;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 28;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S29;
      end
      retro_main_b1_S29: begin
        _address_addr <= 29;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 29;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S30;
      end
      retro_main_b1_S30: begin
        _address_addr <= 30;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 30;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S31;
      end
      retro_main_b1_S31: begin
        _address_addr <= 31;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 31;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S32;
      end
      retro_main_b1_S32: begin
        _address_addr <= 32;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 32;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S33;
      end
      retro_main_b1_S33: begin
        _address_addr <= 33;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 33;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S34;
      end
      retro_main_b1_S34: begin
        _address_addr <= 34;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 34;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S35;
      end
      retro_main_b1_S35: begin
        _address_addr <= 35;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 35;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S36;
      end
      retro_main_b1_S36: begin
        _address_addr <= 36;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 36;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S37;
      end
      retro_main_b1_S37: begin
        _address_addr <= 37;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 37;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S38;
      end
      retro_main_b1_S38: begin
        _address_addr <= 38;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 38;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S39;
      end
      retro_main_b1_S39: begin
        _address_addr <= 39;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 39;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S40;
      end
      retro_main_b1_S40: begin
        _address_addr <= 40;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 40;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S41;
      end
      retro_main_b1_S41: begin
        _address_addr <= 41;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 41;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S42;
      end
      retro_main_b1_S42: begin
        _address_addr <= 42;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 42;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S43;
      end
      retro_main_b1_S43: begin
        _address_addr <= 43;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 43;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S44;
      end
      retro_main_b1_S44: begin
        _address_addr <= 44;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 44;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S45;
      end
      retro_main_b1_S45: begin
        _address_addr <= 45;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 45;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S46;
      end
      retro_main_b1_S46: begin
        _address_addr <= 46;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 46;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S47;
      end
      retro_main_b1_S47: begin
        _address_addr <= 47;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 47;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S48;
      end
      retro_main_b1_S48: begin
        _address_addr <= 48;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 48;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S49;
      end
      retro_main_b1_S49: begin
        _address_addr <= 49;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 49;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S50;
      end
      retro_main_b1_S50: begin
        _address_addr <= 50;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 50;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S51;
      end
      retro_main_b1_S51: begin
        _address_addr <= 51;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 51;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S52;
      end
      retro_main_b1_S52: begin
        _address_addr <= 52;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 52;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S53;
      end
      retro_main_b1_S53: begin
        _address_addr <= 53;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 53;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S54;
      end
      retro_main_b1_S54: begin
        _address_addr <= 54;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 54;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S55;
      end
      retro_main_b1_S55: begin
        _address_addr <= 55;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 55;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S56;
      end
      retro_main_b1_S56: begin
        _address_addr <= 56;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 56;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S57;
      end
      retro_main_b1_S57: begin
        _address_addr <= 57;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 57;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S58;
      end
      retro_main_b1_S58: begin
        _address_addr <= 58;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 58;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S59;
      end
      retro_main_b1_S59: begin
        _address_addr <= 59;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 59;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S60;
      end
      retro_main_b1_S60: begin
        _address_addr <= 60;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 60;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S61;
      end
      retro_main_b1_S61: begin
        _address_addr <= 61;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 61;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S62;
      end
      retro_main_b1_S62: begin
        _address_addr <= 62;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 62;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S63;
      end
      retro_main_b1_S63: begin
        _address_addr <= 63;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 63;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S64;
      end
      retro_main_b1_S64: begin
        _address_addr <= 64;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 64;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S65;
      end
      retro_main_b1_S65: begin
        _address_addr <= 65;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 65;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S66;
      end
      retro_main_b1_S66: begin
        _address_addr <= 66;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 66;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S67;
      end
      retro_main_b1_S67: begin
        _address_addr <= 67;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 67;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S68;
      end
      retro_main_b1_S68: begin
        _address_addr <= 68;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 68;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S69;
      end
      retro_main_b1_S69: begin
        _address_addr <= 69;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 69;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S70;
      end
      retro_main_b1_S70: begin
        _address_addr <= 70;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 70;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S71;
      end
      retro_main_b1_S71: begin
        _address_addr <= 71;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 71;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S72;
      end
      retro_main_b1_S72: begin
        _address_addr <= 72;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 72;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S73;
      end
      retro_main_b1_S73: begin
        _address_addr <= 73;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 73;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S74;
      end
      retro_main_b1_S74: begin
        _address_addr <= 74;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 74;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S75;
      end
      retro_main_b1_S75: begin
        _address_addr <= 75;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 75;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S76;
      end
      retro_main_b1_S76: begin
        _address_addr <= 76;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 76;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S77;
      end
      retro_main_b1_S77: begin
        _address_addr <= 77;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 77;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S78;
      end
      retro_main_b1_S78: begin
        _address_addr <= 78;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 78;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S79;
      end
      retro_main_b1_S79: begin
        _address_addr <= 79;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 79;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S80;
      end
      retro_main_b1_S80: begin
        _address_addr <= 80;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 80;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S81;
      end
      retro_main_b1_S81: begin
        _address_addr <= 81;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 81;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S82;
      end
      retro_main_b1_S82: begin
        _address_addr <= 82;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 82;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S83;
      end
      retro_main_b1_S83: begin
        _address_addr <= 83;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 83;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S84;
      end
      retro_main_b1_S84: begin
        _address_addr <= 84;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 84;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S85;
      end
      retro_main_b1_S85: begin
        _address_addr <= 85;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 85;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S86;
      end
      retro_main_b1_S86: begin
        _address_addr <= 86;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 86;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S87;
      end
      retro_main_b1_S87: begin
        _address_addr <= 87;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 87;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S88;
      end
      retro_main_b1_S88: begin
        _address_addr <= 88;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 88;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S89;
      end
      retro_main_b1_S89: begin
        _address_addr <= 89;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 89;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S90;
      end
      retro_main_b1_S90: begin
        _address_addr <= 90;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 90;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S91;
      end
      retro_main_b1_S91: begin
        _address_addr <= 91;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 91;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S92;
      end
      retro_main_b1_S92: begin
        _address_addr <= 92;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 92;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S93;
      end
      retro_main_b1_S93: begin
        _address_addr <= 93;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 93;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S94;
      end
      retro_main_b1_S94: begin
        _address_addr <= 94;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 94;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S95;
      end
      retro_main_b1_S95: begin
        _address_addr <= 95;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 95;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S96;
      end
      retro_main_b1_S96: begin
        _address_addr <= 96;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 96;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S97;
      end
      retro_main_b1_S97: begin
        _address_addr <= 97;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 97;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S98;
      end
      retro_main_b1_S98: begin
        _address_addr <= 98;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 98;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S99;
      end
      retro_main_b1_S99: begin
        _address_addr <= 99;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 99;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S100;
      end
      retro_main_b1_S100: begin
        _address_addr <= 100;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 100;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S101;
      end
      retro_main_b1_S101: begin
        _address_addr <= 101;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 101;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S102;
      end
      retro_main_b1_S102: begin
        _address_addr <= 102;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 102;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S103;
      end
      retro_main_b1_S103: begin
        _address_addr <= 103;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 103;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S104;
      end
      retro_main_b1_S104: begin
        _address_addr <= 104;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 104;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S105;
      end
      retro_main_b1_S105: begin
        _address_addr <= 105;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 105;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S106;
      end
      retro_main_b1_S106: begin
        _address_addr <= 106;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 106;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S107;
      end
      retro_main_b1_S107: begin
        _address_addr <= 107;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 107;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S108;
      end
      retro_main_b1_S108: begin
        _address_addr <= 108;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 108;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S109;
      end
      retro_main_b1_S109: begin
        _address_addr <= 109;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 109;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S110;
      end
      retro_main_b1_S110: begin
        _address_addr <= 110;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 110;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S111;
      end
      retro_main_b1_S111: begin
        _address_addr <= 111;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 111;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S112;
      end
      retro_main_b1_S112: begin
        _address_addr <= 112;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 112;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S113;
      end
      retro_main_b1_S113: begin
        _address_addr <= 113;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 113;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S114;
      end
      retro_main_b1_S114: begin
        _address_addr <= 114;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 114;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S115;
      end
      retro_main_b1_S115: begin
        _address_addr <= 115;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 115;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S116;
      end
      retro_main_b1_S116: begin
        _address_addr <= 116;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 116;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S117;
      end
      retro_main_b1_S117: begin
        _address_addr <= 117;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 117;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S118;
      end
      retro_main_b1_S118: begin
        _address_addr <= 118;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 118;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S119;
      end
      retro_main_b1_S119: begin
        _address_addr <= 119;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 119;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S120;
      end
      retro_main_b1_S120: begin
        _address_addr <= 120;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 120;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S121;
      end
      retro_main_b1_S121: begin
        _address_addr <= 121;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 121;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S122;
      end
      retro_main_b1_S122: begin
        _address_addr <= 122;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 122;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S123;
      end
      retro_main_b1_S123: begin
        _address_addr <= 123;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 123;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S124;
      end
      retro_main_b1_S124: begin
        _address_addr <= 124;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 124;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S125;
      end
      retro_main_b1_S125: begin
        _address_addr <= 125;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 125;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S126;
      end
      retro_main_b1_S126: begin
        _address_addr <= 126;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 126;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S127;
      end
      retro_main_b1_S127: begin
        _address_addr <= 127;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_addr <= 127;
        _stack_we <= 1;
        _stack_req <= 1;
        _stack_d <= 0;
        retro_main_state <= retro_main_b1_S128;
      end
      retro_main_b1_S128: begin
        _address_addr <= 128;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        _stack_req <= 0;
        retro_main_state <= retro_main_b1_S129;
      end
      retro_main_b1_S129: begin
        _address_addr <= 129;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S130;
      end
      retro_main_b1_S130: begin
        _address_addr <= 130;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S131;
      end
      retro_main_b1_S131: begin
        _address_addr <= 131;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S132;
      end
      retro_main_b1_S132: begin
        _address_addr <= 132;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S133;
      end
      retro_main_b1_S133: begin
        _address_addr <= 133;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S134;
      end
      retro_main_b1_S134: begin
        _address_addr <= 134;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S135;
      end
      retro_main_b1_S135: begin
        _address_addr <= 135;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S136;
      end
      retro_main_b1_S136: begin
        _address_addr <= 136;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S137;
      end
      retro_main_b1_S137: begin
        _address_addr <= 137;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S138;
      end
      retro_main_b1_S138: begin
        _address_addr <= 138;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S139;
      end
      retro_main_b1_S139: begin
        _address_addr <= 139;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S140;
      end
      retro_main_b1_S140: begin
        _address_addr <= 140;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S141;
      end
      retro_main_b1_S141: begin
        _address_addr <= 141;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S142;
      end
      retro_main_b1_S142: begin
        _address_addr <= 142;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S143;
      end
      retro_main_b1_S143: begin
        _address_addr <= 143;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S144;
      end
      retro_main_b1_S144: begin
        _address_addr <= 144;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S145;
      end
      retro_main_b1_S145: begin
        _address_addr <= 145;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S146;
      end
      retro_main_b1_S146: begin
        _address_addr <= 146;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S147;
      end
      retro_main_b1_S147: begin
        _address_addr <= 147;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S148;
      end
      retro_main_b1_S148: begin
        _address_addr <= 148;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S149;
      end
      retro_main_b1_S149: begin
        _address_addr <= 149;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S150;
      end
      retro_main_b1_S150: begin
        _address_addr <= 150;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S151;
      end
      retro_main_b1_S151: begin
        _address_addr <= 151;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S152;
      end
      retro_main_b1_S152: begin
        _address_addr <= 152;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S153;
      end
      retro_main_b1_S153: begin
        _address_addr <= 153;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S154;
      end
      retro_main_b1_S154: begin
        _address_addr <= 154;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S155;
      end
      retro_main_b1_S155: begin
        _address_addr <= 155;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S156;
      end
      retro_main_b1_S156: begin
        _address_addr <= 156;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S157;
      end
      retro_main_b1_S157: begin
        _address_addr <= 157;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S158;
      end
      retro_main_b1_S158: begin
        _address_addr <= 158;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S159;
      end
      retro_main_b1_S159: begin
        _address_addr <= 159;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S160;
      end
      retro_main_b1_S160: begin
        _address_addr <= 160;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S161;
      end
      retro_main_b1_S161: begin
        _address_addr <= 161;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S162;
      end
      retro_main_b1_S162: begin
        _address_addr <= 162;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S163;
      end
      retro_main_b1_S163: begin
        _address_addr <= 163;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S164;
      end
      retro_main_b1_S164: begin
        _address_addr <= 164;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S165;
      end
      retro_main_b1_S165: begin
        _address_addr <= 165;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S166;
      end
      retro_main_b1_S166: begin
        _address_addr <= 166;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S167;
      end
      retro_main_b1_S167: begin
        _address_addr <= 167;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S168;
      end
      retro_main_b1_S168: begin
        _address_addr <= 168;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S169;
      end
      retro_main_b1_S169: begin
        _address_addr <= 169;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S170;
      end
      retro_main_b1_S170: begin
        _address_addr <= 170;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S171;
      end
      retro_main_b1_S171: begin
        _address_addr <= 171;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S172;
      end
      retro_main_b1_S172: begin
        _address_addr <= 172;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S173;
      end
      retro_main_b1_S173: begin
        _address_addr <= 173;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S174;
      end
      retro_main_b1_S174: begin
        _address_addr <= 174;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S175;
      end
      retro_main_b1_S175: begin
        _address_addr <= 175;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S176;
      end
      retro_main_b1_S176: begin
        _address_addr <= 176;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S177;
      end
      retro_main_b1_S177: begin
        _address_addr <= 177;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S178;
      end
      retro_main_b1_S178: begin
        _address_addr <= 178;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S179;
      end
      retro_main_b1_S179: begin
        _address_addr <= 179;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S180;
      end
      retro_main_b1_S180: begin
        _address_addr <= 180;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S181;
      end
      retro_main_b1_S181: begin
        _address_addr <= 181;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S182;
      end
      retro_main_b1_S182: begin
        _address_addr <= 182;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S183;
      end
      retro_main_b1_S183: begin
        _address_addr <= 183;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S184;
      end
      retro_main_b1_S184: begin
        _address_addr <= 184;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S185;
      end
      retro_main_b1_S185: begin
        _address_addr <= 185;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S186;
      end
      retro_main_b1_S186: begin
        _address_addr <= 186;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S187;
      end
      retro_main_b1_S187: begin
        _address_addr <= 187;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S188;
      end
      retro_main_b1_S188: begin
        _address_addr <= 188;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S189;
      end
      retro_main_b1_S189: begin
        _address_addr <= 189;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S190;
      end
      retro_main_b1_S190: begin
        _address_addr <= 190;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S191;
      end
      retro_main_b1_S191: begin
        _address_addr <= 191;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S192;
      end
      retro_main_b1_S192: begin
        _address_addr <= 192;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S193;
      end
      retro_main_b1_S193: begin
        _address_addr <= 193;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S194;
      end
      retro_main_b1_S194: begin
        _address_addr <= 194;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S195;
      end
      retro_main_b1_S195: begin
        _address_addr <= 195;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S196;
      end
      retro_main_b1_S196: begin
        _address_addr <= 196;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S197;
      end
      retro_main_b1_S197: begin
        _address_addr <= 197;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S198;
      end
      retro_main_b1_S198: begin
        _address_addr <= 198;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S199;
      end
      retro_main_b1_S199: begin
        _address_addr <= 199;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S200;
      end
      retro_main_b1_S200: begin
        _address_addr <= 200;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S201;
      end
      retro_main_b1_S201: begin
        _address_addr <= 201;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S202;
      end
      retro_main_b1_S202: begin
        _address_addr <= 202;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S203;
      end
      retro_main_b1_S203: begin
        _address_addr <= 203;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S204;
      end
      retro_main_b1_S204: begin
        _address_addr <= 204;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S205;
      end
      retro_main_b1_S205: begin
        _address_addr <= 205;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S206;
      end
      retro_main_b1_S206: begin
        _address_addr <= 206;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S207;
      end
      retro_main_b1_S207: begin
        _address_addr <= 207;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S208;
      end
      retro_main_b1_S208: begin
        _address_addr <= 208;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S209;
      end
      retro_main_b1_S209: begin
        _address_addr <= 209;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S210;
      end
      retro_main_b1_S210: begin
        _address_addr <= 210;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S211;
      end
      retro_main_b1_S211: begin
        _address_addr <= 211;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S212;
      end
      retro_main_b1_S212: begin
        _address_addr <= 212;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S213;
      end
      retro_main_b1_S213: begin
        _address_addr <= 213;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S214;
      end
      retro_main_b1_S214: begin
        _address_addr <= 214;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S215;
      end
      retro_main_b1_S215: begin
        _address_addr <= 215;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S216;
      end
      retro_main_b1_S216: begin
        _address_addr <= 216;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S217;
      end
      retro_main_b1_S217: begin
        _address_addr <= 217;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S218;
      end
      retro_main_b1_S218: begin
        _address_addr <= 218;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S219;
      end
      retro_main_b1_S219: begin
        _address_addr <= 219;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S220;
      end
      retro_main_b1_S220: begin
        _address_addr <= 220;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S221;
      end
      retro_main_b1_S221: begin
        _address_addr <= 221;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S222;
      end
      retro_main_b1_S222: begin
        _address_addr <= 222;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S223;
      end
      retro_main_b1_S223: begin
        _address_addr <= 223;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S224;
      end
      retro_main_b1_S224: begin
        _address_addr <= 224;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S225;
      end
      retro_main_b1_S225: begin
        _address_addr <= 225;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S226;
      end
      retro_main_b1_S226: begin
        _address_addr <= 226;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S227;
      end
      retro_main_b1_S227: begin
        _address_addr <= 227;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S228;
      end
      retro_main_b1_S228: begin
        _address_addr <= 228;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S229;
      end
      retro_main_b1_S229: begin
        _address_addr <= 229;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S230;
      end
      retro_main_b1_S230: begin
        _address_addr <= 230;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S231;
      end
      retro_main_b1_S231: begin
        _address_addr <= 231;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S232;
      end
      retro_main_b1_S232: begin
        _address_addr <= 232;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S233;
      end
      retro_main_b1_S233: begin
        _address_addr <= 233;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S234;
      end
      retro_main_b1_S234: begin
        _address_addr <= 234;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S235;
      end
      retro_main_b1_S235: begin
        _address_addr <= 235;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S236;
      end
      retro_main_b1_S236: begin
        _address_addr <= 236;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S237;
      end
      retro_main_b1_S237: begin
        _address_addr <= 237;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S238;
      end
      retro_main_b1_S238: begin
        _address_addr <= 238;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S239;
      end
      retro_main_b1_S239: begin
        _address_addr <= 239;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S240;
      end
      retro_main_b1_S240: begin
        _address_addr <= 240;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S241;
      end
      retro_main_b1_S241: begin
        _address_addr <= 241;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S242;
      end
      retro_main_b1_S242: begin
        _address_addr <= 242;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S243;
      end
      retro_main_b1_S243: begin
        _address_addr <= 243;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S244;
      end
      retro_main_b1_S244: begin
        _address_addr <= 244;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S245;
      end
      retro_main_b1_S245: begin
        _address_addr <= 245;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S246;
      end
      retro_main_b1_S246: begin
        _address_addr <= 246;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S247;
      end
      retro_main_b1_S247: begin
        _address_addr <= 247;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S248;
      end
      retro_main_b1_S248: begin
        _address_addr <= 248;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S249;
      end
      retro_main_b1_S249: begin
        _address_addr <= 249;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S250;
      end
      retro_main_b1_S250: begin
        _address_addr <= 250;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S251;
      end
      retro_main_b1_S251: begin
        _address_addr <= 251;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S252;
      end
      retro_main_b1_S252: begin
        _address_addr <= 252;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S253;
      end
      retro_main_b1_S253: begin
        _address_addr <= 253;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S254;
      end
      retro_main_b1_S254: begin
        _address_addr <= 254;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S255;
      end
      retro_main_b1_S255: begin
        _address_addr <= 255;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S256;
      end
      retro_main_b1_S256: begin
        _address_addr <= 256;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S257;
      end
      retro_main_b1_S257: begin
        _address_addr <= 257;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S258;
      end
      retro_main_b1_S258: begin
        _address_addr <= 258;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S259;
      end
      retro_main_b1_S259: begin
        _address_addr <= 259;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S260;
      end
      retro_main_b1_S260: begin
        _address_addr <= 260;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S261;
      end
      retro_main_b1_S261: begin
        _address_addr <= 261;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S262;
      end
      retro_main_b1_S262: begin
        _address_addr <= 262;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S263;
      end
      retro_main_b1_S263: begin
        _address_addr <= 263;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S264;
      end
      retro_main_b1_S264: begin
        _address_addr <= 264;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S265;
      end
      retro_main_b1_S265: begin
        _address_addr <= 265;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S266;
      end
      retro_main_b1_S266: begin
        _address_addr <= 266;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S267;
      end
      retro_main_b1_S267: begin
        _address_addr <= 267;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S268;
      end
      retro_main_b1_S268: begin
        _address_addr <= 268;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S269;
      end
      retro_main_b1_S269: begin
        _address_addr <= 269;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S270;
      end
      retro_main_b1_S270: begin
        _address_addr <= 270;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S271;
      end
      retro_main_b1_S271: begin
        _address_addr <= 271;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S272;
      end
      retro_main_b1_S272: begin
        _address_addr <= 272;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S273;
      end
      retro_main_b1_S273: begin
        _address_addr <= 273;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S274;
      end
      retro_main_b1_S274: begin
        _address_addr <= 274;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S275;
      end
      retro_main_b1_S275: begin
        _address_addr <= 275;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S276;
      end
      retro_main_b1_S276: begin
        _address_addr <= 276;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S277;
      end
      retro_main_b1_S277: begin
        _address_addr <= 277;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S278;
      end
      retro_main_b1_S278: begin
        _address_addr <= 278;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S279;
      end
      retro_main_b1_S279: begin
        _address_addr <= 279;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S280;
      end
      retro_main_b1_S280: begin
        _address_addr <= 280;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S281;
      end
      retro_main_b1_S281: begin
        _address_addr <= 281;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S282;
      end
      retro_main_b1_S282: begin
        _address_addr <= 282;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S283;
      end
      retro_main_b1_S283: begin
        _address_addr <= 283;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S284;
      end
      retro_main_b1_S284: begin
        _address_addr <= 284;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S285;
      end
      retro_main_b1_S285: begin
        _address_addr <= 285;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S286;
      end
      retro_main_b1_S286: begin
        _address_addr <= 286;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S287;
      end
      retro_main_b1_S287: begin
        _address_addr <= 287;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S288;
      end
      retro_main_b1_S288: begin
        _address_addr <= 288;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S289;
      end
      retro_main_b1_S289: begin
        _address_addr <= 289;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S290;
      end
      retro_main_b1_S290: begin
        _address_addr <= 290;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S291;
      end
      retro_main_b1_S291: begin
        _address_addr <= 291;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S292;
      end
      retro_main_b1_S292: begin
        _address_addr <= 292;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S293;
      end
      retro_main_b1_S293: begin
        _address_addr <= 293;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S294;
      end
      retro_main_b1_S294: begin
        _address_addr <= 294;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S295;
      end
      retro_main_b1_S295: begin
        _address_addr <= 295;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S296;
      end
      retro_main_b1_S296: begin
        _address_addr <= 296;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S297;
      end
      retro_main_b1_S297: begin
        _address_addr <= 297;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S298;
      end
      retro_main_b1_S298: begin
        _address_addr <= 298;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S299;
      end
      retro_main_b1_S299: begin
        _address_addr <= 299;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S300;
      end
      retro_main_b1_S300: begin
        _address_addr <= 300;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S301;
      end
      retro_main_b1_S301: begin
        _address_addr <= 301;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S302;
      end
      retro_main_b1_S302: begin
        _address_addr <= 302;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S303;
      end
      retro_main_b1_S303: begin
        _address_addr <= 303;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S304;
      end
      retro_main_b1_S304: begin
        _address_addr <= 304;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S305;
      end
      retro_main_b1_S305: begin
        _address_addr <= 305;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S306;
      end
      retro_main_b1_S306: begin
        _address_addr <= 306;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S307;
      end
      retro_main_b1_S307: begin
        _address_addr <= 307;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S308;
      end
      retro_main_b1_S308: begin
        _address_addr <= 308;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S309;
      end
      retro_main_b1_S309: begin
        _address_addr <= 309;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S310;
      end
      retro_main_b1_S310: begin
        _address_addr <= 310;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S311;
      end
      retro_main_b1_S311: begin
        _address_addr <= 311;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S312;
      end
      retro_main_b1_S312: begin
        _address_addr <= 312;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S313;
      end
      retro_main_b1_S313: begin
        _address_addr <= 313;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S314;
      end
      retro_main_b1_S314: begin
        _address_addr <= 314;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S315;
      end
      retro_main_b1_S315: begin
        _address_addr <= 315;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S316;
      end
      retro_main_b1_S316: begin
        _address_addr <= 316;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S317;
      end
      retro_main_b1_S317: begin
        _address_addr <= 317;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S318;
      end
      retro_main_b1_S318: begin
        _address_addr <= 318;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S319;
      end
      retro_main_b1_S319: begin
        _address_addr <= 319;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S320;
      end
      retro_main_b1_S320: begin
        _address_addr <= 320;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S321;
      end
      retro_main_b1_S321: begin
        _address_addr <= 321;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S322;
      end
      retro_main_b1_S322: begin
        _address_addr <= 322;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S323;
      end
      retro_main_b1_S323: begin
        _address_addr <= 323;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S324;
      end
      retro_main_b1_S324: begin
        _address_addr <= 324;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S325;
      end
      retro_main_b1_S325: begin
        _address_addr <= 325;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S326;
      end
      retro_main_b1_S326: begin
        _address_addr <= 326;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S327;
      end
      retro_main_b1_S327: begin
        _address_addr <= 327;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S328;
      end
      retro_main_b1_S328: begin
        _address_addr <= 328;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S329;
      end
      retro_main_b1_S329: begin
        _address_addr <= 329;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S330;
      end
      retro_main_b1_S330: begin
        _address_addr <= 330;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S331;
      end
      retro_main_b1_S331: begin
        _address_addr <= 331;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S332;
      end
      retro_main_b1_S332: begin
        _address_addr <= 332;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S333;
      end
      retro_main_b1_S333: begin
        _address_addr <= 333;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S334;
      end
      retro_main_b1_S334: begin
        _address_addr <= 334;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S335;
      end
      retro_main_b1_S335: begin
        _address_addr <= 335;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S336;
      end
      retro_main_b1_S336: begin
        _address_addr <= 336;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S337;
      end
      retro_main_b1_S337: begin
        _address_addr <= 337;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S338;
      end
      retro_main_b1_S338: begin
        _address_addr <= 338;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S339;
      end
      retro_main_b1_S339: begin
        _address_addr <= 339;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S340;
      end
      retro_main_b1_S340: begin
        _address_addr <= 340;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S341;
      end
      retro_main_b1_S341: begin
        _address_addr <= 341;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S342;
      end
      retro_main_b1_S342: begin
        _address_addr <= 342;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S343;
      end
      retro_main_b1_S343: begin
        _address_addr <= 343;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S344;
      end
      retro_main_b1_S344: begin
        _address_addr <= 344;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S345;
      end
      retro_main_b1_S345: begin
        _address_addr <= 345;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S346;
      end
      retro_main_b1_S346: begin
        _address_addr <= 346;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S347;
      end
      retro_main_b1_S347: begin
        _address_addr <= 347;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S348;
      end
      retro_main_b1_S348: begin
        _address_addr <= 348;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S349;
      end
      retro_main_b1_S349: begin
        _address_addr <= 349;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S350;
      end
      retro_main_b1_S350: begin
        _address_addr <= 350;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S351;
      end
      retro_main_b1_S351: begin
        _address_addr <= 351;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S352;
      end
      retro_main_b1_S352: begin
        _address_addr <= 352;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S353;
      end
      retro_main_b1_S353: begin
        _address_addr <= 353;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S354;
      end
      retro_main_b1_S354: begin
        _address_addr <= 354;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S355;
      end
      retro_main_b1_S355: begin
        _address_addr <= 355;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S356;
      end
      retro_main_b1_S356: begin
        _address_addr <= 356;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S357;
      end
      retro_main_b1_S357: begin
        _address_addr <= 357;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S358;
      end
      retro_main_b1_S358: begin
        _address_addr <= 358;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S359;
      end
      retro_main_b1_S359: begin
        _address_addr <= 359;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S360;
      end
      retro_main_b1_S360: begin
        _address_addr <= 360;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S361;
      end
      retro_main_b1_S361: begin
        _address_addr <= 361;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S362;
      end
      retro_main_b1_S362: begin
        _address_addr <= 362;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S363;
      end
      retro_main_b1_S363: begin
        _address_addr <= 363;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S364;
      end
      retro_main_b1_S364: begin
        _address_addr <= 364;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S365;
      end
      retro_main_b1_S365: begin
        _address_addr <= 365;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S366;
      end
      retro_main_b1_S366: begin
        _address_addr <= 366;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S367;
      end
      retro_main_b1_S367: begin
        _address_addr <= 367;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S368;
      end
      retro_main_b1_S368: begin
        _address_addr <= 368;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S369;
      end
      retro_main_b1_S369: begin
        _address_addr <= 369;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S370;
      end
      retro_main_b1_S370: begin
        _address_addr <= 370;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S371;
      end
      retro_main_b1_S371: begin
        _address_addr <= 371;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S372;
      end
      retro_main_b1_S372: begin
        _address_addr <= 372;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S373;
      end
      retro_main_b1_S373: begin
        _address_addr <= 373;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S374;
      end
      retro_main_b1_S374: begin
        _address_addr <= 374;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S375;
      end
      retro_main_b1_S375: begin
        _address_addr <= 375;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S376;
      end
      retro_main_b1_S376: begin
        _address_addr <= 376;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S377;
      end
      retro_main_b1_S377: begin
        _address_addr <= 377;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S378;
      end
      retro_main_b1_S378: begin
        _address_addr <= 378;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S379;
      end
      retro_main_b1_S379: begin
        _address_addr <= 379;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S380;
      end
      retro_main_b1_S380: begin
        _address_addr <= 380;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S381;
      end
      retro_main_b1_S381: begin
        _address_addr <= 381;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S382;
      end
      retro_main_b1_S382: begin
        _address_addr <= 382;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S383;
      end
      retro_main_b1_S383: begin
        _address_addr <= 383;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S384;
      end
      retro_main_b1_S384: begin
        _address_addr <= 384;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S385;
      end
      retro_main_b1_S385: begin
        _address_addr <= 385;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S386;
      end
      retro_main_b1_S386: begin
        _address_addr <= 386;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S387;
      end
      retro_main_b1_S387: begin
        _address_addr <= 387;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S388;
      end
      retro_main_b1_S388: begin
        _address_addr <= 388;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S389;
      end
      retro_main_b1_S389: begin
        _address_addr <= 389;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S390;
      end
      retro_main_b1_S390: begin
        _address_addr <= 390;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S391;
      end
      retro_main_b1_S391: begin
        _address_addr <= 391;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S392;
      end
      retro_main_b1_S392: begin
        _address_addr <= 392;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S393;
      end
      retro_main_b1_S393: begin
        _address_addr <= 393;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S394;
      end
      retro_main_b1_S394: begin
        _address_addr <= 394;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S395;
      end
      retro_main_b1_S395: begin
        _address_addr <= 395;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S396;
      end
      retro_main_b1_S396: begin
        _address_addr <= 396;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S397;
      end
      retro_main_b1_S397: begin
        _address_addr <= 397;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S398;
      end
      retro_main_b1_S398: begin
        _address_addr <= 398;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S399;
      end
      retro_main_b1_S399: begin
        _address_addr <= 399;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S400;
      end
      retro_main_b1_S400: begin
        _address_addr <= 400;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S401;
      end
      retro_main_b1_S401: begin
        _address_addr <= 401;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S402;
      end
      retro_main_b1_S402: begin
        _address_addr <= 402;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S403;
      end
      retro_main_b1_S403: begin
        _address_addr <= 403;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S404;
      end
      retro_main_b1_S404: begin
        _address_addr <= 404;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S405;
      end
      retro_main_b1_S405: begin
        _address_addr <= 405;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S406;
      end
      retro_main_b1_S406: begin
        _address_addr <= 406;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S407;
      end
      retro_main_b1_S407: begin
        _address_addr <= 407;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S408;
      end
      retro_main_b1_S408: begin
        _address_addr <= 408;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S409;
      end
      retro_main_b1_S409: begin
        _address_addr <= 409;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S410;
      end
      retro_main_b1_S410: begin
        _address_addr <= 410;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S411;
      end
      retro_main_b1_S411: begin
        _address_addr <= 411;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S412;
      end
      retro_main_b1_S412: begin
        _address_addr <= 412;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S413;
      end
      retro_main_b1_S413: begin
        _address_addr <= 413;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S414;
      end
      retro_main_b1_S414: begin
        _address_addr <= 414;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S415;
      end
      retro_main_b1_S415: begin
        _address_addr <= 415;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S416;
      end
      retro_main_b1_S416: begin
        _address_addr <= 416;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S417;
      end
      retro_main_b1_S417: begin
        _address_addr <= 417;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S418;
      end
      retro_main_b1_S418: begin
        _address_addr <= 418;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S419;
      end
      retro_main_b1_S419: begin
        _address_addr <= 419;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S420;
      end
      retro_main_b1_S420: begin
        _address_addr <= 420;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S421;
      end
      retro_main_b1_S421: begin
        _address_addr <= 421;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S422;
      end
      retro_main_b1_S422: begin
        _address_addr <= 422;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S423;
      end
      retro_main_b1_S423: begin
        _address_addr <= 423;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S424;
      end
      retro_main_b1_S424: begin
        _address_addr <= 424;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S425;
      end
      retro_main_b1_S425: begin
        _address_addr <= 425;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S426;
      end
      retro_main_b1_S426: begin
        _address_addr <= 426;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S427;
      end
      retro_main_b1_S427: begin
        _address_addr <= 427;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S428;
      end
      retro_main_b1_S428: begin
        _address_addr <= 428;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S429;
      end
      retro_main_b1_S429: begin
        _address_addr <= 429;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S430;
      end
      retro_main_b1_S430: begin
        _address_addr <= 430;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S431;
      end
      retro_main_b1_S431: begin
        _address_addr <= 431;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S432;
      end
      retro_main_b1_S432: begin
        _address_addr <= 432;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S433;
      end
      retro_main_b1_S433: begin
        _address_addr <= 433;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S434;
      end
      retro_main_b1_S434: begin
        _address_addr <= 434;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S435;
      end
      retro_main_b1_S435: begin
        _address_addr <= 435;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S436;
      end
      retro_main_b1_S436: begin
        _address_addr <= 436;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S437;
      end
      retro_main_b1_S437: begin
        _address_addr <= 437;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S438;
      end
      retro_main_b1_S438: begin
        _address_addr <= 438;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S439;
      end
      retro_main_b1_S439: begin
        _address_addr <= 439;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S440;
      end
      retro_main_b1_S440: begin
        _address_addr <= 440;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S441;
      end
      retro_main_b1_S441: begin
        _address_addr <= 441;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S442;
      end
      retro_main_b1_S442: begin
        _address_addr <= 442;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S443;
      end
      retro_main_b1_S443: begin
        _address_addr <= 443;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S444;
      end
      retro_main_b1_S444: begin
        _address_addr <= 444;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S445;
      end
      retro_main_b1_S445: begin
        _address_addr <= 445;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S446;
      end
      retro_main_b1_S446: begin
        _address_addr <= 446;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S447;
      end
      retro_main_b1_S447: begin
        _address_addr <= 447;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S448;
      end
      retro_main_b1_S448: begin
        _address_addr <= 448;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S449;
      end
      retro_main_b1_S449: begin
        _address_addr <= 449;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S450;
      end
      retro_main_b1_S450: begin
        _address_addr <= 450;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S451;
      end
      retro_main_b1_S451: begin
        _address_addr <= 451;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S452;
      end
      retro_main_b1_S452: begin
        _address_addr <= 452;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S453;
      end
      retro_main_b1_S453: begin
        _address_addr <= 453;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S454;
      end
      retro_main_b1_S454: begin
        _address_addr <= 454;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S455;
      end
      retro_main_b1_S455: begin
        _address_addr <= 455;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S456;
      end
      retro_main_b1_S456: begin
        _address_addr <= 456;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S457;
      end
      retro_main_b1_S457: begin
        _address_addr <= 457;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S458;
      end
      retro_main_b1_S458: begin
        _address_addr <= 458;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S459;
      end
      retro_main_b1_S459: begin
        _address_addr <= 459;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S460;
      end
      retro_main_b1_S460: begin
        _address_addr <= 460;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S461;
      end
      retro_main_b1_S461: begin
        _address_addr <= 461;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S462;
      end
      retro_main_b1_S462: begin
        _address_addr <= 462;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S463;
      end
      retro_main_b1_S463: begin
        _address_addr <= 463;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S464;
      end
      retro_main_b1_S464: begin
        _address_addr <= 464;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S465;
      end
      retro_main_b1_S465: begin
        _address_addr <= 465;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S466;
      end
      retro_main_b1_S466: begin
        _address_addr <= 466;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S467;
      end
      retro_main_b1_S467: begin
        _address_addr <= 467;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S468;
      end
      retro_main_b1_S468: begin
        _address_addr <= 468;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S469;
      end
      retro_main_b1_S469: begin
        _address_addr <= 469;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S470;
      end
      retro_main_b1_S470: begin
        _address_addr <= 470;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S471;
      end
      retro_main_b1_S471: begin
        _address_addr <= 471;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S472;
      end
      retro_main_b1_S472: begin
        _address_addr <= 472;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S473;
      end
      retro_main_b1_S473: begin
        _address_addr <= 473;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S474;
      end
      retro_main_b1_S474: begin
        _address_addr <= 474;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S475;
      end
      retro_main_b1_S475: begin
        _address_addr <= 475;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S476;
      end
      retro_main_b1_S476: begin
        _address_addr <= 476;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S477;
      end
      retro_main_b1_S477: begin
        _address_addr <= 477;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S478;
      end
      retro_main_b1_S478: begin
        _address_addr <= 478;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S479;
      end
      retro_main_b1_S479: begin
        _address_addr <= 479;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S480;
      end
      retro_main_b1_S480: begin
        _address_addr <= 480;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S481;
      end
      retro_main_b1_S481: begin
        _address_addr <= 481;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S482;
      end
      retro_main_b1_S482: begin
        _address_addr <= 482;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S483;
      end
      retro_main_b1_S483: begin
        _address_addr <= 483;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S484;
      end
      retro_main_b1_S484: begin
        _address_addr <= 484;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S485;
      end
      retro_main_b1_S485: begin
        _address_addr <= 485;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S486;
      end
      retro_main_b1_S486: begin
        _address_addr <= 486;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S487;
      end
      retro_main_b1_S487: begin
        _address_addr <= 487;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S488;
      end
      retro_main_b1_S488: begin
        _address_addr <= 488;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S489;
      end
      retro_main_b1_S489: begin
        _address_addr <= 489;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S490;
      end
      retro_main_b1_S490: begin
        _address_addr <= 490;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S491;
      end
      retro_main_b1_S491: begin
        _address_addr <= 491;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S492;
      end
      retro_main_b1_S492: begin
        _address_addr <= 492;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S493;
      end
      retro_main_b1_S493: begin
        _address_addr <= 493;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S494;
      end
      retro_main_b1_S494: begin
        _address_addr <= 494;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S495;
      end
      retro_main_b1_S495: begin
        _address_addr <= 495;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S496;
      end
      retro_main_b1_S496: begin
        _address_addr <= 496;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S497;
      end
      retro_main_b1_S497: begin
        _address_addr <= 497;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S498;
      end
      retro_main_b1_S498: begin
        _address_addr <= 498;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S499;
      end
      retro_main_b1_S499: begin
        _address_addr <= 499;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S500;
      end
      retro_main_b1_S500: begin
        _address_addr <= 500;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S501;
      end
      retro_main_b1_S501: begin
        _address_addr <= 501;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S502;
      end
      retro_main_b1_S502: begin
        _address_addr <= 502;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S503;
      end
      retro_main_b1_S503: begin
        _address_addr <= 503;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S504;
      end
      retro_main_b1_S504: begin
        _address_addr <= 504;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S505;
      end
      retro_main_b1_S505: begin
        _address_addr <= 505;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S506;
      end
      retro_main_b1_S506: begin
        _address_addr <= 506;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S507;
      end
      retro_main_b1_S507: begin
        _address_addr <= 507;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S508;
      end
      retro_main_b1_S508: begin
        _address_addr <= 508;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S509;
      end
      retro_main_b1_S509: begin
        _address_addr <= 509;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S510;
      end
      retro_main_b1_S510: begin
        _address_addr <= 510;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S511;
      end
      retro_main_b1_S511: begin
        _address_addr <= 511;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S512;
      end
      retro_main_b1_S512: begin
        _address_addr <= 512;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S513;
      end
      retro_main_b1_S513: begin
        _address_addr <= 513;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S514;
      end
      retro_main_b1_S514: begin
        _address_addr <= 514;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S515;
      end
      retro_main_b1_S515: begin
        _address_addr <= 515;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S516;
      end
      retro_main_b1_S516: begin
        _address_addr <= 516;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S517;
      end
      retro_main_b1_S517: begin
        _address_addr <= 517;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S518;
      end
      retro_main_b1_S518: begin
        _address_addr <= 518;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S519;
      end
      retro_main_b1_S519: begin
        _address_addr <= 519;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S520;
      end
      retro_main_b1_S520: begin
        _address_addr <= 520;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S521;
      end
      retro_main_b1_S521: begin
        _address_addr <= 521;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S522;
      end
      retro_main_b1_S522: begin
        _address_addr <= 522;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S523;
      end
      retro_main_b1_S523: begin
        _address_addr <= 523;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S524;
      end
      retro_main_b1_S524: begin
        _address_addr <= 524;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S525;
      end
      retro_main_b1_S525: begin
        _address_addr <= 525;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S526;
      end
      retro_main_b1_S526: begin
        _address_addr <= 526;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S527;
      end
      retro_main_b1_S527: begin
        _address_addr <= 527;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S528;
      end
      retro_main_b1_S528: begin
        _address_addr <= 528;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S529;
      end
      retro_main_b1_S529: begin
        _address_addr <= 529;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S530;
      end
      retro_main_b1_S530: begin
        _address_addr <= 530;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S531;
      end
      retro_main_b1_S531: begin
        _address_addr <= 531;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S532;
      end
      retro_main_b1_S532: begin
        _address_addr <= 532;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S533;
      end
      retro_main_b1_S533: begin
        _address_addr <= 533;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S534;
      end
      retro_main_b1_S534: begin
        _address_addr <= 534;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S535;
      end
      retro_main_b1_S535: begin
        _address_addr <= 535;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S536;
      end
      retro_main_b1_S536: begin
        _address_addr <= 536;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S537;
      end
      retro_main_b1_S537: begin
        _address_addr <= 537;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S538;
      end
      retro_main_b1_S538: begin
        _address_addr <= 538;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S539;
      end
      retro_main_b1_S539: begin
        _address_addr <= 539;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S540;
      end
      retro_main_b1_S540: begin
        _address_addr <= 540;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S541;
      end
      retro_main_b1_S541: begin
        _address_addr <= 541;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S542;
      end
      retro_main_b1_S542: begin
        _address_addr <= 542;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S543;
      end
      retro_main_b1_S543: begin
        _address_addr <= 543;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S544;
      end
      retro_main_b1_S544: begin
        _address_addr <= 544;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S545;
      end
      retro_main_b1_S545: begin
        _address_addr <= 545;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S546;
      end
      retro_main_b1_S546: begin
        _address_addr <= 546;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S547;
      end
      retro_main_b1_S547: begin
        _address_addr <= 547;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S548;
      end
      retro_main_b1_S548: begin
        _address_addr <= 548;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S549;
      end
      retro_main_b1_S549: begin
        _address_addr <= 549;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S550;
      end
      retro_main_b1_S550: begin
        _address_addr <= 550;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S551;
      end
      retro_main_b1_S551: begin
        _address_addr <= 551;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S552;
      end
      retro_main_b1_S552: begin
        _address_addr <= 552;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S553;
      end
      retro_main_b1_S553: begin
        _address_addr <= 553;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S554;
      end
      retro_main_b1_S554: begin
        _address_addr <= 554;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S555;
      end
      retro_main_b1_S555: begin
        _address_addr <= 555;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S556;
      end
      retro_main_b1_S556: begin
        _address_addr <= 556;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S557;
      end
      retro_main_b1_S557: begin
        _address_addr <= 557;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S558;
      end
      retro_main_b1_S558: begin
        _address_addr <= 558;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S559;
      end
      retro_main_b1_S559: begin
        _address_addr <= 559;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S560;
      end
      retro_main_b1_S560: begin
        _address_addr <= 560;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S561;
      end
      retro_main_b1_S561: begin
        _address_addr <= 561;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S562;
      end
      retro_main_b1_S562: begin
        _address_addr <= 562;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S563;
      end
      retro_main_b1_S563: begin
        _address_addr <= 563;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S564;
      end
      retro_main_b1_S564: begin
        _address_addr <= 564;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S565;
      end
      retro_main_b1_S565: begin
        _address_addr <= 565;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S566;
      end
      retro_main_b1_S566: begin
        _address_addr <= 566;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S567;
      end
      retro_main_b1_S567: begin
        _address_addr <= 567;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S568;
      end
      retro_main_b1_S568: begin
        _address_addr <= 568;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S569;
      end
      retro_main_b1_S569: begin
        _address_addr <= 569;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S570;
      end
      retro_main_b1_S570: begin
        _address_addr <= 570;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S571;
      end
      retro_main_b1_S571: begin
        _address_addr <= 571;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S572;
      end
      retro_main_b1_S572: begin
        _address_addr <= 572;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S573;
      end
      retro_main_b1_S573: begin
        _address_addr <= 573;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S574;
      end
      retro_main_b1_S574: begin
        _address_addr <= 574;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S575;
      end
      retro_main_b1_S575: begin
        _address_addr <= 575;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S576;
      end
      retro_main_b1_S576: begin
        _address_addr <= 576;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S577;
      end
      retro_main_b1_S577: begin
        _address_addr <= 577;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S578;
      end
      retro_main_b1_S578: begin
        _address_addr <= 578;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S579;
      end
      retro_main_b1_S579: begin
        _address_addr <= 579;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S580;
      end
      retro_main_b1_S580: begin
        _address_addr <= 580;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S581;
      end
      retro_main_b1_S581: begin
        _address_addr <= 581;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S582;
      end
      retro_main_b1_S582: begin
        _address_addr <= 582;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S583;
      end
      retro_main_b1_S583: begin
        _address_addr <= 583;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S584;
      end
      retro_main_b1_S584: begin
        _address_addr <= 584;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S585;
      end
      retro_main_b1_S585: begin
        _address_addr <= 585;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S586;
      end
      retro_main_b1_S586: begin
        _address_addr <= 586;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S587;
      end
      retro_main_b1_S587: begin
        _address_addr <= 587;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S588;
      end
      retro_main_b1_S588: begin
        _address_addr <= 588;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S589;
      end
      retro_main_b1_S589: begin
        _address_addr <= 589;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S590;
      end
      retro_main_b1_S590: begin
        _address_addr <= 590;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S591;
      end
      retro_main_b1_S591: begin
        _address_addr <= 591;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S592;
      end
      retro_main_b1_S592: begin
        _address_addr <= 592;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S593;
      end
      retro_main_b1_S593: begin
        _address_addr <= 593;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S594;
      end
      retro_main_b1_S594: begin
        _address_addr <= 594;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S595;
      end
      retro_main_b1_S595: begin
        _address_addr <= 595;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S596;
      end
      retro_main_b1_S596: begin
        _address_addr <= 596;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S597;
      end
      retro_main_b1_S597: begin
        _address_addr <= 597;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S598;
      end
      retro_main_b1_S598: begin
        _address_addr <= 598;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S599;
      end
      retro_main_b1_S599: begin
        _address_addr <= 599;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S600;
      end
      retro_main_b1_S600: begin
        _address_addr <= 600;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S601;
      end
      retro_main_b1_S601: begin
        _address_addr <= 601;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S602;
      end
      retro_main_b1_S602: begin
        _address_addr <= 602;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S603;
      end
      retro_main_b1_S603: begin
        _address_addr <= 603;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S604;
      end
      retro_main_b1_S604: begin
        _address_addr <= 604;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S605;
      end
      retro_main_b1_S605: begin
        _address_addr <= 605;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S606;
      end
      retro_main_b1_S606: begin
        _address_addr <= 606;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S607;
      end
      retro_main_b1_S607: begin
        _address_addr <= 607;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S608;
      end
      retro_main_b1_S608: begin
        _address_addr <= 608;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S609;
      end
      retro_main_b1_S609: begin
        _address_addr <= 609;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S610;
      end
      retro_main_b1_S610: begin
        _address_addr <= 610;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S611;
      end
      retro_main_b1_S611: begin
        _address_addr <= 611;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S612;
      end
      retro_main_b1_S612: begin
        _address_addr <= 612;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S613;
      end
      retro_main_b1_S613: begin
        _address_addr <= 613;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S614;
      end
      retro_main_b1_S614: begin
        _address_addr <= 614;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S615;
      end
      retro_main_b1_S615: begin
        _address_addr <= 615;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S616;
      end
      retro_main_b1_S616: begin
        _address_addr <= 616;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S617;
      end
      retro_main_b1_S617: begin
        _address_addr <= 617;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S618;
      end
      retro_main_b1_S618: begin
        _address_addr <= 618;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S619;
      end
      retro_main_b1_S619: begin
        _address_addr <= 619;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S620;
      end
      retro_main_b1_S620: begin
        _address_addr <= 620;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S621;
      end
      retro_main_b1_S621: begin
        _address_addr <= 621;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S622;
      end
      retro_main_b1_S622: begin
        _address_addr <= 622;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S623;
      end
      retro_main_b1_S623: begin
        _address_addr <= 623;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S624;
      end
      retro_main_b1_S624: begin
        _address_addr <= 624;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S625;
      end
      retro_main_b1_S625: begin
        _address_addr <= 625;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S626;
      end
      retro_main_b1_S626: begin
        _address_addr <= 626;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S627;
      end
      retro_main_b1_S627: begin
        _address_addr <= 627;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S628;
      end
      retro_main_b1_S628: begin
        _address_addr <= 628;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S629;
      end
      retro_main_b1_S629: begin
        _address_addr <= 629;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S630;
      end
      retro_main_b1_S630: begin
        _address_addr <= 630;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S631;
      end
      retro_main_b1_S631: begin
        _address_addr <= 631;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S632;
      end
      retro_main_b1_S632: begin
        _address_addr <= 632;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S633;
      end
      retro_main_b1_S633: begin
        _address_addr <= 633;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S634;
      end
      retro_main_b1_S634: begin
        _address_addr <= 634;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S635;
      end
      retro_main_b1_S635: begin
        _address_addr <= 635;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S636;
      end
      retro_main_b1_S636: begin
        _address_addr <= 636;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S637;
      end
      retro_main_b1_S637: begin
        _address_addr <= 637;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S638;
      end
      retro_main_b1_S638: begin
        _address_addr <= 638;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S639;
      end
      retro_main_b1_S639: begin
        _address_addr <= 639;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S640;
      end
      retro_main_b1_S640: begin
        _address_addr <= 640;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S641;
      end
      retro_main_b1_S641: begin
        _address_addr <= 641;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S642;
      end
      retro_main_b1_S642: begin
        _address_addr <= 642;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S643;
      end
      retro_main_b1_S643: begin
        _address_addr <= 643;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S644;
      end
      retro_main_b1_S644: begin
        _address_addr <= 644;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S645;
      end
      retro_main_b1_S645: begin
        _address_addr <= 645;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S646;
      end
      retro_main_b1_S646: begin
        _address_addr <= 646;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S647;
      end
      retro_main_b1_S647: begin
        _address_addr <= 647;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S648;
      end
      retro_main_b1_S648: begin
        _address_addr <= 648;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S649;
      end
      retro_main_b1_S649: begin
        _address_addr <= 649;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S650;
      end
      retro_main_b1_S650: begin
        _address_addr <= 650;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S651;
      end
      retro_main_b1_S651: begin
        _address_addr <= 651;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S652;
      end
      retro_main_b1_S652: begin
        _address_addr <= 652;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S653;
      end
      retro_main_b1_S653: begin
        _address_addr <= 653;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S654;
      end
      retro_main_b1_S654: begin
        _address_addr <= 654;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S655;
      end
      retro_main_b1_S655: begin
        _address_addr <= 655;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S656;
      end
      retro_main_b1_S656: begin
        _address_addr <= 656;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S657;
      end
      retro_main_b1_S657: begin
        _address_addr <= 657;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S658;
      end
      retro_main_b1_S658: begin
        _address_addr <= 658;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S659;
      end
      retro_main_b1_S659: begin
        _address_addr <= 659;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S660;
      end
      retro_main_b1_S660: begin
        _address_addr <= 660;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S661;
      end
      retro_main_b1_S661: begin
        _address_addr <= 661;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S662;
      end
      retro_main_b1_S662: begin
        _address_addr <= 662;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S663;
      end
      retro_main_b1_S663: begin
        _address_addr <= 663;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S664;
      end
      retro_main_b1_S664: begin
        _address_addr <= 664;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S665;
      end
      retro_main_b1_S665: begin
        _address_addr <= 665;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S666;
      end
      retro_main_b1_S666: begin
        _address_addr <= 666;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S667;
      end
      retro_main_b1_S667: begin
        _address_addr <= 667;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S668;
      end
      retro_main_b1_S668: begin
        _address_addr <= 668;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S669;
      end
      retro_main_b1_S669: begin
        _address_addr <= 669;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S670;
      end
      retro_main_b1_S670: begin
        _address_addr <= 670;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S671;
      end
      retro_main_b1_S671: begin
        _address_addr <= 671;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S672;
      end
      retro_main_b1_S672: begin
        _address_addr <= 672;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S673;
      end
      retro_main_b1_S673: begin
        _address_addr <= 673;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S674;
      end
      retro_main_b1_S674: begin
        _address_addr <= 674;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S675;
      end
      retro_main_b1_S675: begin
        _address_addr <= 675;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S676;
      end
      retro_main_b1_S676: begin
        _address_addr <= 676;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S677;
      end
      retro_main_b1_S677: begin
        _address_addr <= 677;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S678;
      end
      retro_main_b1_S678: begin
        _address_addr <= 678;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S679;
      end
      retro_main_b1_S679: begin
        _address_addr <= 679;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S680;
      end
      retro_main_b1_S680: begin
        _address_addr <= 680;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S681;
      end
      retro_main_b1_S681: begin
        _address_addr <= 681;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S682;
      end
      retro_main_b1_S682: begin
        _address_addr <= 682;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S683;
      end
      retro_main_b1_S683: begin
        _address_addr <= 683;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S684;
      end
      retro_main_b1_S684: begin
        _address_addr <= 684;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S685;
      end
      retro_main_b1_S685: begin
        _address_addr <= 685;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S686;
      end
      retro_main_b1_S686: begin
        _address_addr <= 686;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S687;
      end
      retro_main_b1_S687: begin
        _address_addr <= 687;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S688;
      end
      retro_main_b1_S688: begin
        _address_addr <= 688;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S689;
      end
      retro_main_b1_S689: begin
        _address_addr <= 689;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S690;
      end
      retro_main_b1_S690: begin
        _address_addr <= 690;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S691;
      end
      retro_main_b1_S691: begin
        _address_addr <= 691;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S692;
      end
      retro_main_b1_S692: begin
        _address_addr <= 692;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S693;
      end
      retro_main_b1_S693: begin
        _address_addr <= 693;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S694;
      end
      retro_main_b1_S694: begin
        _address_addr <= 694;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S695;
      end
      retro_main_b1_S695: begin
        _address_addr <= 695;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S696;
      end
      retro_main_b1_S696: begin
        _address_addr <= 696;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S697;
      end
      retro_main_b1_S697: begin
        _address_addr <= 697;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S698;
      end
      retro_main_b1_S698: begin
        _address_addr <= 698;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S699;
      end
      retro_main_b1_S699: begin
        _address_addr <= 699;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S700;
      end
      retro_main_b1_S700: begin
        _address_addr <= 700;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S701;
      end
      retro_main_b1_S701: begin
        _address_addr <= 701;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S702;
      end
      retro_main_b1_S702: begin
        _address_addr <= 702;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S703;
      end
      retro_main_b1_S703: begin
        _address_addr <= 703;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S704;
      end
      retro_main_b1_S704: begin
        _address_addr <= 704;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S705;
      end
      retro_main_b1_S705: begin
        _address_addr <= 705;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S706;
      end
      retro_main_b1_S706: begin
        _address_addr <= 706;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S707;
      end
      retro_main_b1_S707: begin
        _address_addr <= 707;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S708;
      end
      retro_main_b1_S708: begin
        _address_addr <= 708;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S709;
      end
      retro_main_b1_S709: begin
        _address_addr <= 709;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S710;
      end
      retro_main_b1_S710: begin
        _address_addr <= 710;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S711;
      end
      retro_main_b1_S711: begin
        _address_addr <= 711;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S712;
      end
      retro_main_b1_S712: begin
        _address_addr <= 712;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S713;
      end
      retro_main_b1_S713: begin
        _address_addr <= 713;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S714;
      end
      retro_main_b1_S714: begin
        _address_addr <= 714;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S715;
      end
      retro_main_b1_S715: begin
        _address_addr <= 715;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S716;
      end
      retro_main_b1_S716: begin
        _address_addr <= 716;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S717;
      end
      retro_main_b1_S717: begin
        _address_addr <= 717;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S718;
      end
      retro_main_b1_S718: begin
        _address_addr <= 718;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S719;
      end
      retro_main_b1_S719: begin
        _address_addr <= 719;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S720;
      end
      retro_main_b1_S720: begin
        _address_addr <= 720;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S721;
      end
      retro_main_b1_S721: begin
        _address_addr <= 721;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S722;
      end
      retro_main_b1_S722: begin
        _address_addr <= 722;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S723;
      end
      retro_main_b1_S723: begin
        _address_addr <= 723;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S724;
      end
      retro_main_b1_S724: begin
        _address_addr <= 724;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S725;
      end
      retro_main_b1_S725: begin
        _address_addr <= 725;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S726;
      end
      retro_main_b1_S726: begin
        _address_addr <= 726;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S727;
      end
      retro_main_b1_S727: begin
        _address_addr <= 727;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S728;
      end
      retro_main_b1_S728: begin
        _address_addr <= 728;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S729;
      end
      retro_main_b1_S729: begin
        _address_addr <= 729;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S730;
      end
      retro_main_b1_S730: begin
        _address_addr <= 730;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S731;
      end
      retro_main_b1_S731: begin
        _address_addr <= 731;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S732;
      end
      retro_main_b1_S732: begin
        _address_addr <= 732;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S733;
      end
      retro_main_b1_S733: begin
        _address_addr <= 733;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S734;
      end
      retro_main_b1_S734: begin
        _address_addr <= 734;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S735;
      end
      retro_main_b1_S735: begin
        _address_addr <= 735;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S736;
      end
      retro_main_b1_S736: begin
        _address_addr <= 736;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S737;
      end
      retro_main_b1_S737: begin
        _address_addr <= 737;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S738;
      end
      retro_main_b1_S738: begin
        _address_addr <= 738;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S739;
      end
      retro_main_b1_S739: begin
        _address_addr <= 739;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S740;
      end
      retro_main_b1_S740: begin
        _address_addr <= 740;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S741;
      end
      retro_main_b1_S741: begin
        _address_addr <= 741;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S742;
      end
      retro_main_b1_S742: begin
        _address_addr <= 742;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S743;
      end
      retro_main_b1_S743: begin
        _address_addr <= 743;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S744;
      end
      retro_main_b1_S744: begin
        _address_addr <= 744;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S745;
      end
      retro_main_b1_S745: begin
        _address_addr <= 745;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S746;
      end
      retro_main_b1_S746: begin
        _address_addr <= 746;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S747;
      end
      retro_main_b1_S747: begin
        _address_addr <= 747;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S748;
      end
      retro_main_b1_S748: begin
        _address_addr <= 748;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S749;
      end
      retro_main_b1_S749: begin
        _address_addr <= 749;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S750;
      end
      retro_main_b1_S750: begin
        _address_addr <= 750;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S751;
      end
      retro_main_b1_S751: begin
        _address_addr <= 751;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S752;
      end
      retro_main_b1_S752: begin
        _address_addr <= 752;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S753;
      end
      retro_main_b1_S753: begin
        _address_addr <= 753;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S754;
      end
      retro_main_b1_S754: begin
        _address_addr <= 754;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S755;
      end
      retro_main_b1_S755: begin
        _address_addr <= 755;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S756;
      end
      retro_main_b1_S756: begin
        _address_addr <= 756;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S757;
      end
      retro_main_b1_S757: begin
        _address_addr <= 757;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S758;
      end
      retro_main_b1_S758: begin
        _address_addr <= 758;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S759;
      end
      retro_main_b1_S759: begin
        _address_addr <= 759;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S760;
      end
      retro_main_b1_S760: begin
        _address_addr <= 760;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S761;
      end
      retro_main_b1_S761: begin
        _address_addr <= 761;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S762;
      end
      retro_main_b1_S762: begin
        _address_addr <= 762;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S763;
      end
      retro_main_b1_S763: begin
        _address_addr <= 763;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S764;
      end
      retro_main_b1_S764: begin
        _address_addr <= 764;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S765;
      end
      retro_main_b1_S765: begin
        _address_addr <= 765;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S766;
      end
      retro_main_b1_S766: begin
        _address_addr <= 766;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S767;
      end
      retro_main_b1_S767: begin
        _address_addr <= 767;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S768;
      end
      retro_main_b1_S768: begin
        _address_addr <= 768;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S769;
      end
      retro_main_b1_S769: begin
        _address_addr <= 769;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S770;
      end
      retro_main_b1_S770: begin
        _address_addr <= 770;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S771;
      end
      retro_main_b1_S771: begin
        _address_addr <= 771;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S772;
      end
      retro_main_b1_S772: begin
        _address_addr <= 772;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S773;
      end
      retro_main_b1_S773: begin
        _address_addr <= 773;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S774;
      end
      retro_main_b1_S774: begin
        _address_addr <= 774;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S775;
      end
      retro_main_b1_S775: begin
        _address_addr <= 775;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S776;
      end
      retro_main_b1_S776: begin
        _address_addr <= 776;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S777;
      end
      retro_main_b1_S777: begin
        _address_addr <= 777;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S778;
      end
      retro_main_b1_S778: begin
        _address_addr <= 778;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S779;
      end
      retro_main_b1_S779: begin
        _address_addr <= 779;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S780;
      end
      retro_main_b1_S780: begin
        _address_addr <= 780;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S781;
      end
      retro_main_b1_S781: begin
        _address_addr <= 781;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S782;
      end
      retro_main_b1_S782: begin
        _address_addr <= 782;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S783;
      end
      retro_main_b1_S783: begin
        _address_addr <= 783;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S784;
      end
      retro_main_b1_S784: begin
        _address_addr <= 784;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S785;
      end
      retro_main_b1_S785: begin
        _address_addr <= 785;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S786;
      end
      retro_main_b1_S786: begin
        _address_addr <= 786;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S787;
      end
      retro_main_b1_S787: begin
        _address_addr <= 787;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S788;
      end
      retro_main_b1_S788: begin
        _address_addr <= 788;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S789;
      end
      retro_main_b1_S789: begin
        _address_addr <= 789;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S790;
      end
      retro_main_b1_S790: begin
        _address_addr <= 790;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S791;
      end
      retro_main_b1_S791: begin
        _address_addr <= 791;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S792;
      end
      retro_main_b1_S792: begin
        _address_addr <= 792;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S793;
      end
      retro_main_b1_S793: begin
        _address_addr <= 793;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S794;
      end
      retro_main_b1_S794: begin
        _address_addr <= 794;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S795;
      end
      retro_main_b1_S795: begin
        _address_addr <= 795;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S796;
      end
      retro_main_b1_S796: begin
        _address_addr <= 796;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S797;
      end
      retro_main_b1_S797: begin
        _address_addr <= 797;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S798;
      end
      retro_main_b1_S798: begin
        _address_addr <= 798;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S799;
      end
      retro_main_b1_S799: begin
        _address_addr <= 799;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S800;
      end
      retro_main_b1_S800: begin
        _address_addr <= 800;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S801;
      end
      retro_main_b1_S801: begin
        _address_addr <= 801;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S802;
      end
      retro_main_b1_S802: begin
        _address_addr <= 802;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S803;
      end
      retro_main_b1_S803: begin
        _address_addr <= 803;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S804;
      end
      retro_main_b1_S804: begin
        _address_addr <= 804;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S805;
      end
      retro_main_b1_S805: begin
        _address_addr <= 805;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S806;
      end
      retro_main_b1_S806: begin
        _address_addr <= 806;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S807;
      end
      retro_main_b1_S807: begin
        _address_addr <= 807;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S808;
      end
      retro_main_b1_S808: begin
        _address_addr <= 808;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S809;
      end
      retro_main_b1_S809: begin
        _address_addr <= 809;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S810;
      end
      retro_main_b1_S810: begin
        _address_addr <= 810;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S811;
      end
      retro_main_b1_S811: begin
        _address_addr <= 811;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S812;
      end
      retro_main_b1_S812: begin
        _address_addr <= 812;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S813;
      end
      retro_main_b1_S813: begin
        _address_addr <= 813;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S814;
      end
      retro_main_b1_S814: begin
        _address_addr <= 814;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S815;
      end
      retro_main_b1_S815: begin
        _address_addr <= 815;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S816;
      end
      retro_main_b1_S816: begin
        _address_addr <= 816;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S817;
      end
      retro_main_b1_S817: begin
        _address_addr <= 817;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S818;
      end
      retro_main_b1_S818: begin
        _address_addr <= 818;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S819;
      end
      retro_main_b1_S819: begin
        _address_addr <= 819;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S820;
      end
      retro_main_b1_S820: begin
        _address_addr <= 820;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S821;
      end
      retro_main_b1_S821: begin
        _address_addr <= 821;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S822;
      end
      retro_main_b1_S822: begin
        _address_addr <= 822;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S823;
      end
      retro_main_b1_S823: begin
        _address_addr <= 823;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S824;
      end
      retro_main_b1_S824: begin
        _address_addr <= 824;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S825;
      end
      retro_main_b1_S825: begin
        _address_addr <= 825;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S826;
      end
      retro_main_b1_S826: begin
        _address_addr <= 826;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S827;
      end
      retro_main_b1_S827: begin
        _address_addr <= 827;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S828;
      end
      retro_main_b1_S828: begin
        _address_addr <= 828;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S829;
      end
      retro_main_b1_S829: begin
        _address_addr <= 829;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S830;
      end
      retro_main_b1_S830: begin
        _address_addr <= 830;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S831;
      end
      retro_main_b1_S831: begin
        _address_addr <= 831;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S832;
      end
      retro_main_b1_S832: begin
        _address_addr <= 832;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S833;
      end
      retro_main_b1_S833: begin
        _address_addr <= 833;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S834;
      end
      retro_main_b1_S834: begin
        _address_addr <= 834;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S835;
      end
      retro_main_b1_S835: begin
        _address_addr <= 835;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S836;
      end
      retro_main_b1_S836: begin
        _address_addr <= 836;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S837;
      end
      retro_main_b1_S837: begin
        _address_addr <= 837;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S838;
      end
      retro_main_b1_S838: begin
        _address_addr <= 838;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S839;
      end
      retro_main_b1_S839: begin
        _address_addr <= 839;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S840;
      end
      retro_main_b1_S840: begin
        _address_addr <= 840;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S841;
      end
      retro_main_b1_S841: begin
        _address_addr <= 841;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S842;
      end
      retro_main_b1_S842: begin
        _address_addr <= 842;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S843;
      end
      retro_main_b1_S843: begin
        _address_addr <= 843;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S844;
      end
      retro_main_b1_S844: begin
        _address_addr <= 844;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S845;
      end
      retro_main_b1_S845: begin
        _address_addr <= 845;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S846;
      end
      retro_main_b1_S846: begin
        _address_addr <= 846;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S847;
      end
      retro_main_b1_S847: begin
        _address_addr <= 847;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S848;
      end
      retro_main_b1_S848: begin
        _address_addr <= 848;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S849;
      end
      retro_main_b1_S849: begin
        _address_addr <= 849;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S850;
      end
      retro_main_b1_S850: begin
        _address_addr <= 850;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S851;
      end
      retro_main_b1_S851: begin
        _address_addr <= 851;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S852;
      end
      retro_main_b1_S852: begin
        _address_addr <= 852;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S853;
      end
      retro_main_b1_S853: begin
        _address_addr <= 853;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S854;
      end
      retro_main_b1_S854: begin
        _address_addr <= 854;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S855;
      end
      retro_main_b1_S855: begin
        _address_addr <= 855;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S856;
      end
      retro_main_b1_S856: begin
        _address_addr <= 856;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S857;
      end
      retro_main_b1_S857: begin
        _address_addr <= 857;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S858;
      end
      retro_main_b1_S858: begin
        _address_addr <= 858;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S859;
      end
      retro_main_b1_S859: begin
        _address_addr <= 859;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S860;
      end
      retro_main_b1_S860: begin
        _address_addr <= 860;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S861;
      end
      retro_main_b1_S861: begin
        _address_addr <= 861;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S862;
      end
      retro_main_b1_S862: begin
        _address_addr <= 862;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S863;
      end
      retro_main_b1_S863: begin
        _address_addr <= 863;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S864;
      end
      retro_main_b1_S864: begin
        _address_addr <= 864;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S865;
      end
      retro_main_b1_S865: begin
        _address_addr <= 865;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S866;
      end
      retro_main_b1_S866: begin
        _address_addr <= 866;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S867;
      end
      retro_main_b1_S867: begin
        _address_addr <= 867;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S868;
      end
      retro_main_b1_S868: begin
        _address_addr <= 868;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S869;
      end
      retro_main_b1_S869: begin
        _address_addr <= 869;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S870;
      end
      retro_main_b1_S870: begin
        _address_addr <= 870;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S871;
      end
      retro_main_b1_S871: begin
        _address_addr <= 871;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S872;
      end
      retro_main_b1_S872: begin
        _address_addr <= 872;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S873;
      end
      retro_main_b1_S873: begin
        _address_addr <= 873;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S874;
      end
      retro_main_b1_S874: begin
        _address_addr <= 874;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S875;
      end
      retro_main_b1_S875: begin
        _address_addr <= 875;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S876;
      end
      retro_main_b1_S876: begin
        _address_addr <= 876;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S877;
      end
      retro_main_b1_S877: begin
        _address_addr <= 877;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S878;
      end
      retro_main_b1_S878: begin
        _address_addr <= 878;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S879;
      end
      retro_main_b1_S879: begin
        _address_addr <= 879;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S880;
      end
      retro_main_b1_S880: begin
        _address_addr <= 880;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S881;
      end
      retro_main_b1_S881: begin
        _address_addr <= 881;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S882;
      end
      retro_main_b1_S882: begin
        _address_addr <= 882;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S883;
      end
      retro_main_b1_S883: begin
        _address_addr <= 883;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S884;
      end
      retro_main_b1_S884: begin
        _address_addr <= 884;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S885;
      end
      retro_main_b1_S885: begin
        _address_addr <= 885;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S886;
      end
      retro_main_b1_S886: begin
        _address_addr <= 886;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S887;
      end
      retro_main_b1_S887: begin
        _address_addr <= 887;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S888;
      end
      retro_main_b1_S888: begin
        _address_addr <= 888;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S889;
      end
      retro_main_b1_S889: begin
        _address_addr <= 889;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S890;
      end
      retro_main_b1_S890: begin
        _address_addr <= 890;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S891;
      end
      retro_main_b1_S891: begin
        _address_addr <= 891;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S892;
      end
      retro_main_b1_S892: begin
        _address_addr <= 892;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S893;
      end
      retro_main_b1_S893: begin
        _address_addr <= 893;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S894;
      end
      retro_main_b1_S894: begin
        _address_addr <= 894;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S895;
      end
      retro_main_b1_S895: begin
        _address_addr <= 895;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S896;
      end
      retro_main_b1_S896: begin
        _address_addr <= 896;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S897;
      end
      retro_main_b1_S897: begin
        _address_addr <= 897;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S898;
      end
      retro_main_b1_S898: begin
        _address_addr <= 898;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S899;
      end
      retro_main_b1_S899: begin
        _address_addr <= 899;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S900;
      end
      retro_main_b1_S900: begin
        _address_addr <= 900;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S901;
      end
      retro_main_b1_S901: begin
        _address_addr <= 901;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S902;
      end
      retro_main_b1_S902: begin
        _address_addr <= 902;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S903;
      end
      retro_main_b1_S903: begin
        _address_addr <= 903;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S904;
      end
      retro_main_b1_S904: begin
        _address_addr <= 904;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S905;
      end
      retro_main_b1_S905: begin
        _address_addr <= 905;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S906;
      end
      retro_main_b1_S906: begin
        _address_addr <= 906;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S907;
      end
      retro_main_b1_S907: begin
        _address_addr <= 907;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S908;
      end
      retro_main_b1_S908: begin
        _address_addr <= 908;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S909;
      end
      retro_main_b1_S909: begin
        _address_addr <= 909;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S910;
      end
      retro_main_b1_S910: begin
        _address_addr <= 910;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S911;
      end
      retro_main_b1_S911: begin
        _address_addr <= 911;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S912;
      end
      retro_main_b1_S912: begin
        _address_addr <= 912;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S913;
      end
      retro_main_b1_S913: begin
        _address_addr <= 913;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S914;
      end
      retro_main_b1_S914: begin
        _address_addr <= 914;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S915;
      end
      retro_main_b1_S915: begin
        _address_addr <= 915;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S916;
      end
      retro_main_b1_S916: begin
        _address_addr <= 916;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S917;
      end
      retro_main_b1_S917: begin
        _address_addr <= 917;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S918;
      end
      retro_main_b1_S918: begin
        _address_addr <= 918;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S919;
      end
      retro_main_b1_S919: begin
        _address_addr <= 919;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S920;
      end
      retro_main_b1_S920: begin
        _address_addr <= 920;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S921;
      end
      retro_main_b1_S921: begin
        _address_addr <= 921;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S922;
      end
      retro_main_b1_S922: begin
        _address_addr <= 922;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S923;
      end
      retro_main_b1_S923: begin
        _address_addr <= 923;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S924;
      end
      retro_main_b1_S924: begin
        _address_addr <= 924;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S925;
      end
      retro_main_b1_S925: begin
        _address_addr <= 925;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S926;
      end
      retro_main_b1_S926: begin
        _address_addr <= 926;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S927;
      end
      retro_main_b1_S927: begin
        _address_addr <= 927;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S928;
      end
      retro_main_b1_S928: begin
        _address_addr <= 928;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S929;
      end
      retro_main_b1_S929: begin
        _address_addr <= 929;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S930;
      end
      retro_main_b1_S930: begin
        _address_addr <= 930;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S931;
      end
      retro_main_b1_S931: begin
        _address_addr <= 931;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S932;
      end
      retro_main_b1_S932: begin
        _address_addr <= 932;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S933;
      end
      retro_main_b1_S933: begin
        _address_addr <= 933;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S934;
      end
      retro_main_b1_S934: begin
        _address_addr <= 934;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S935;
      end
      retro_main_b1_S935: begin
        _address_addr <= 935;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S936;
      end
      retro_main_b1_S936: begin
        _address_addr <= 936;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S937;
      end
      retro_main_b1_S937: begin
        _address_addr <= 937;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S938;
      end
      retro_main_b1_S938: begin
        _address_addr <= 938;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S939;
      end
      retro_main_b1_S939: begin
        _address_addr <= 939;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S940;
      end
      retro_main_b1_S940: begin
        _address_addr <= 940;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S941;
      end
      retro_main_b1_S941: begin
        _address_addr <= 941;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S942;
      end
      retro_main_b1_S942: begin
        _address_addr <= 942;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S943;
      end
      retro_main_b1_S943: begin
        _address_addr <= 943;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S944;
      end
      retro_main_b1_S944: begin
        _address_addr <= 944;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S945;
      end
      retro_main_b1_S945: begin
        _address_addr <= 945;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S946;
      end
      retro_main_b1_S946: begin
        _address_addr <= 946;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S947;
      end
      retro_main_b1_S947: begin
        _address_addr <= 947;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S948;
      end
      retro_main_b1_S948: begin
        _address_addr <= 948;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S949;
      end
      retro_main_b1_S949: begin
        _address_addr <= 949;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S950;
      end
      retro_main_b1_S950: begin
        _address_addr <= 950;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S951;
      end
      retro_main_b1_S951: begin
        _address_addr <= 951;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S952;
      end
      retro_main_b1_S952: begin
        _address_addr <= 952;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S953;
      end
      retro_main_b1_S953: begin
        _address_addr <= 953;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S954;
      end
      retro_main_b1_S954: begin
        _address_addr <= 954;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S955;
      end
      retro_main_b1_S955: begin
        _address_addr <= 955;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S956;
      end
      retro_main_b1_S956: begin
        _address_addr <= 956;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S957;
      end
      retro_main_b1_S957: begin
        _address_addr <= 957;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S958;
      end
      retro_main_b1_S958: begin
        _address_addr <= 958;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S959;
      end
      retro_main_b1_S959: begin
        _address_addr <= 959;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S960;
      end
      retro_main_b1_S960: begin
        _address_addr <= 960;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S961;
      end
      retro_main_b1_S961: begin
        _address_addr <= 961;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S962;
      end
      retro_main_b1_S962: begin
        _address_addr <= 962;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S963;
      end
      retro_main_b1_S963: begin
        _address_addr <= 963;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S964;
      end
      retro_main_b1_S964: begin
        _address_addr <= 964;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S965;
      end
      retro_main_b1_S965: begin
        _address_addr <= 965;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S966;
      end
      retro_main_b1_S966: begin
        _address_addr <= 966;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S967;
      end
      retro_main_b1_S967: begin
        _address_addr <= 967;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S968;
      end
      retro_main_b1_S968: begin
        _address_addr <= 968;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S969;
      end
      retro_main_b1_S969: begin
        _address_addr <= 969;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S970;
      end
      retro_main_b1_S970: begin
        _address_addr <= 970;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S971;
      end
      retro_main_b1_S971: begin
        _address_addr <= 971;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S972;
      end
      retro_main_b1_S972: begin
        _address_addr <= 972;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S973;
      end
      retro_main_b1_S973: begin
        _address_addr <= 973;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S974;
      end
      retro_main_b1_S974: begin
        _address_addr <= 974;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S975;
      end
      retro_main_b1_S975: begin
        _address_addr <= 975;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S976;
      end
      retro_main_b1_S976: begin
        _address_addr <= 976;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S977;
      end
      retro_main_b1_S977: begin
        _address_addr <= 977;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S978;
      end
      retro_main_b1_S978: begin
        _address_addr <= 978;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S979;
      end
      retro_main_b1_S979: begin
        _address_addr <= 979;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S980;
      end
      retro_main_b1_S980: begin
        _address_addr <= 980;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S981;
      end
      retro_main_b1_S981: begin
        _address_addr <= 981;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S982;
      end
      retro_main_b1_S982: begin
        _address_addr <= 982;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S983;
      end
      retro_main_b1_S983: begin
        _address_addr <= 983;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S984;
      end
      retro_main_b1_S984: begin
        _address_addr <= 984;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S985;
      end
      retro_main_b1_S985: begin
        _address_addr <= 985;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S986;
      end
      retro_main_b1_S986: begin
        _address_addr <= 986;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S987;
      end
      retro_main_b1_S987: begin
        _address_addr <= 987;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S988;
      end
      retro_main_b1_S988: begin
        _address_addr <= 988;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S989;
      end
      retro_main_b1_S989: begin
        _address_addr <= 989;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S990;
      end
      retro_main_b1_S990: begin
        _address_addr <= 990;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S991;
      end
      retro_main_b1_S991: begin
        _address_addr <= 991;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S992;
      end
      retro_main_b1_S992: begin
        _address_addr <= 992;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S993;
      end
      retro_main_b1_S993: begin
        _address_addr <= 993;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S994;
      end
      retro_main_b1_S994: begin
        _address_addr <= 994;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S995;
      end
      retro_main_b1_S995: begin
        _address_addr <= 995;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S996;
      end
      retro_main_b1_S996: begin
        _address_addr <= 996;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S997;
      end
      retro_main_b1_S997: begin
        _address_addr <= 997;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S998;
      end
      retro_main_b1_S998: begin
        _address_addr <= 998;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S999;
      end
      retro_main_b1_S999: begin
        _address_addr <= 999;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S1000;
      end
      retro_main_b1_S1000: begin
        _address_addr <= 1000;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S1001;
      end
      retro_main_b1_S1001: begin
        _address_addr <= 1001;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S1002;
      end
      retro_main_b1_S1002: begin
        _address_addr <= 1002;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S1003;
      end
      retro_main_b1_S1003: begin
        _address_addr <= 1003;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S1004;
      end
      retro_main_b1_S1004: begin
        _address_addr <= 1004;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S1005;
      end
      retro_main_b1_S1005: begin
        _address_addr <= 1005;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S1006;
      end
      retro_main_b1_S1006: begin
        _address_addr <= 1006;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S1007;
      end
      retro_main_b1_S1007: begin
        _address_addr <= 1007;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S1008;
      end
      retro_main_b1_S1008: begin
        _address_addr <= 1008;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S1009;
      end
      retro_main_b1_S1009: begin
        _address_addr <= 1009;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S1010;
      end
      retro_main_b1_S1010: begin
        _address_addr <= 1010;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S1011;
      end
      retro_main_b1_S1011: begin
        _address_addr <= 1011;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S1012;
      end
      retro_main_b1_S1012: begin
        _address_addr <= 1012;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S1013;
      end
      retro_main_b1_S1013: begin
        _address_addr <= 1013;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S1014;
      end
      retro_main_b1_S1014: begin
        _address_addr <= 1014;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S1015;
      end
      retro_main_b1_S1015: begin
        _address_addr <= 1015;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S1016;
      end
      retro_main_b1_S1016: begin
        _address_addr <= 1016;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S1017;
      end
      retro_main_b1_S1017: begin
        _address_addr <= 1017;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S1018;
      end
      retro_main_b1_S1018: begin
        _address_addr <= 1018;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S1019;
      end
      retro_main_b1_S1019: begin
        _address_addr <= 1019;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S1020;
      end
      retro_main_b1_S1020: begin
        _address_addr <= 1020;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S1021;
      end
      retro_main_b1_S1021: begin
        _address_addr <= 1021;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S1022;
      end
      retro_main_b1_S1022: begin
        _address_addr <= 1022;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S1023;
      end
      retro_main_b1_S1023: begin
        _address_addr <= 1023;
        _address_we <= 1;
        _address_req <= 1;
        _address_d <= 0;
        retro_main_state <= retro_main_b1_S1024;
      end
      retro_main_b1_S1024: begin
        _address_req <= 0;
        retro_main_state <= retro_main_L1_while2_S0;
      end
      retro_main_L1_while2_S0: begin
        /* c914 <= (ip2 < 16384); */
        if (c914) begin
          io_ports_addr <= 8;
          io_ports_we <= 1;
          io_ports_req <= 1;
          io_ports_d <= ip2;
          memory_addr <= ip2;
          memory_we <= 0;
          memory_req <= 1;
          retro_main_state <= retro_main_L1_whilebody3_S1;
        end else begin
          retro_main_valid <= 1;
          if (retro_main_accept == 1) begin
            retro_main_state <= retro_main_b1_INIT;
          end
        end
      end
      retro_main_L1_whilebody3_S1: begin
        io_ports_req <= 0;
        /*wait for output of memory*/
        retro_main_state <= retro_main_L1_whilebody3_S2;
      end
      retro_main_L1_whilebody3_S2: begin
        opcode3 <= memory_q;
        memory_req <= 0;
        retro_main_state <= retro_main_L1_whilebody3_S3;
      end
      retro_main_L1_whilebody3_S3: begin
        io_ports_addr <= 9;
        io_ports_we <= 1;
        io_ports_req <= 1;
        io_ports_d <= opcode3;
        /* c915 <= (opcode3 <= 30); */
        retro_main_state <= retro_main_L1_whilebody3_S4;
      end
      retro_main_L1_whilebody3_S4: begin
        io_ports_req <= 0;
        if (c915) begin
          /* c916 <= (opcode3 == 0); */
          /* c917 <= (opcode3 == 1); */
          /* c918 <= (opcode3 == 2); */
          /* c919 <= (opcode3 == 3); */
          /* c920 <= (opcode3 == 4); */
          /* c921 <= (opcode3 == 5); */
          /* c922 <= (opcode3 == 6); */
          /* c923 <= (opcode3 == 7); */
          /* c924 <= (opcode3 == 8); */
          /* c925 <= (opcode3 == 9); */
          /* c926 <= (opcode3 == 10); */
          /* c927 <= (opcode3 == 11); */
          /* c928 <= (opcode3 == 12); */
          /* c929 <= (opcode3 == 13); */
          /* c930 <= (opcode3 == 14); */
          /* c931 <= (opcode3 == 15); */
          /* c932 <= (opcode3 == 16); */
          /* c933 <= (opcode3 == 17); */
          /* c934 <= (opcode3 == 18); */
          /* c935 <= (opcode3 == 19); */
          /* c936 <= (opcode3 == 20); */
          /* c937 <= (opcode3 == 21); */
          /* c938 <= (opcode3 == 22); */
          /* c939 <= (opcode3 == 23); */
          /* c940 <= (opcode3 == 24); */
          /* c941 <= (opcode3 == 25); */
          /* c942 <= (opcode3 == 26); */
          /* c943 <= (opcode3 == 27); */
          /* c944 <= (opcode3 == 28); */
          /* c945 <= (opcode3 == 29); */
          /* c946 <= (opcode3 == 30); */
          /* c2856 <= (c914 && c915); */
          /* c2157 <= (c914 && c915); */
          /* c1106 <= (!c916 && c917); */
          /* c1107 <= ((!c916 && !c917) && c918); */
          /* c1108 <= (((!c916 && !c917) && !c918) && c919); */
          /* c1109 <= ((((!c916 && !c917) && !c918) && !c919) && c920); */
          /* c1110 <= (((((!c916 && !c917) && !c918) && !c919) && !c920) && c921); */
          /* c1111 <= ((((((!c916 && !c917) && !c918) && !c919) && !c920) && !c921) && c922); */
          /* c1112 <= (((((((!c916 && !c917) && !c918) && !c919) && !c920) && !c921) && !c922) && c923); */
          /* c1113 <= ((((((((!c916 && !c917) && !c918) && !c919) && !c920) && !c921) && !c922) && !c923) && c924); */
          /* c1114 <= (((((((((!c916 && !c917) && !c918) && !c919) && !c920) && !c921) && !c922) && !c923) && !c924) && c925); */
          /* c1115 <= ((((((((((!c916 && !c917) && !c918) && !c919) && !c920) && !c921) && !c922) && !c923) && !c924) && !c925) && c926); */
          /* c1116 <= (((((((((((!c916 && !c917) && !c918) && !c919) && !c920) && !c921) && !c922) && !c923) && !c924) && !c925) && !c926) && c927); */
          /* c1117 <= ((((((((((((!c916 && !c917) && !c918) && !c919) && !c920) && !c921) && !c922) && !c923) && !c924) && !c925) && !c926) && !c927) && c928); */
          /* c1118 <= (((((((((((((!c916 && !c917) && !c918) && !c919) && !c920) && !c921) && !c922) && !c923) && !c924) && !c925) && !c926) && !c927) && !c928) && c929); */
          /* c1119 <= ((((((((((((((!c916 && !c917) && !c918) && !c919) && !c920) && !c921) && !c922) && !c923) && !c924) && !c925) && !c926) && !c927) && !c928) && !c929) && c930); */
          /* c1120 <= (((((((((((((((!c916 && !c917) && !c918) && !c919) && !c920) && !c921) && !c922) && !c923) && !c924) && !c925) && !c926) && !c927) && !c928) && !c929) && !c930) && c931); */
          /* c1121 <= ((((((((((((((((!c916 && !c917) && !c918) && !c919) && !c920) && !c921) && !c922) && !c923) && !c924) && !c925) && !c926) && !c927) && !c928) && !c929) && !c930) && !c931) && c932); */
          /* c1122 <= (((((((((((((((((!c916 && !c917) && !c918) && !c919) && !c920) && !c921) && !c922) && !c923) && !c924) && !c925) && !c926) && !c927) && !c928) && !c929) && !c930) && !c931) && !c932) && c933); */
          /* c1123 <= ((((((((((((((((((!c916 && !c917) && !c918) && !c919) && !c920) && !c921) && !c922) && !c923) && !c924) && !c925) && !c926) && !c927) && !c928) && !c929) && !c930) && !c931) && !c932) && !c933) && c934); */
          /* c1124 <= (((((((((((((((((((!c916 && !c917) && !c918) && !c919) && !c920) && !c921) && !c922) && !c923) && !c924) && !c925) && !c926) && !c927) && !c928) && !c929) && !c930) && !c931) && !c932) && !c933) && !c934) && c935); */
          /* c1125 <= ((((((((((((((((((((!c916 && !c917) && !c918) && !c919) && !c920) && !c921) && !c922) && !c923) && !c924) && !c925) && !c926) && !c927) && !c928) && !c929) && !c930) && !c931) && !c932) && !c933) && !c934) && !c935) && c936); */
          /* c1126 <= (((((((((((((((((((((!c916 && !c917) && !c918) && !c919) && !c920) && !c921) && !c922) && !c923) && !c924) && !c925) && !c926) && !c927) && !c928) && !c929) && !c930) && !c931) && !c932) && !c933) && !c934) && !c935) && !c936) && c937); */
          /* c1127 <= ((((((((((((((((((((((!c916 && !c917) && !c918) && !c919) && !c920) && !c921) && !c922) && !c923) && !c924) && !c925) && !c926) && !c927) && !c928) && !c929) && !c930) && !c931) && !c932) && !c933) && !c934) && !c935) && !c936) && !c937) && c938); */
          /* c1128 <= (((((((((((((((((((((((!c916 && !c917) && !c918) && !c919) && !c920) && !c921) && !c922) && !c923) && !c924) && !c925) && !c926) && !c927) && !c928) && !c929) && !c930) && !c931) && !c932) && !c933) && !c934) && !c935) && !c936) && !c937) && !c938) && c939); */
          /* c1129 <= ((((((((((((((((((((((((!c916 && !c917) && !c918) && !c919) && !c920) && !c921) && !c922) && !c923) && !c924) && !c925) && !c926) && !c927) && !c928) && !c929) && !c930) && !c931) && !c932) && !c933) && !c934) && !c935) && !c936) && !c937) && !c938) && !c939) && c940); */
          /* c1130 <= (((((((((((((((((((((((((!c916 && !c917) && !c918) && !c919) && !c920) && !c921) && !c922) && !c923) && !c924) && !c925) && !c926) && !c927) && !c928) && !c929) && !c930) && !c931) && !c932) && !c933) && !c934) && !c935) && !c936) && !c937) && !c938) && !c939) && !c940) && c941); */
          /* c1131 <= ((((((((((((((((((((((((((!c916 && !c917) && !c918) && !c919) && !c920) && !c921) && !c922) && !c923) && !c924) && !c925) && !c926) && !c927) && !c928) && !c929) && !c930) && !c931) && !c932) && !c933) && !c934) && !c935) && !c936) && !c937) && !c938) && !c939) && !c940) && !c941) && c942); */
          /* c1132 <= (((((((((((((((((((((((((((!c916 && !c917) && !c918) && !c919) && !c920) && !c921) && !c922) && !c923) && !c924) && !c925) && !c926) && !c927) && !c928) && !c929) && !c930) && !c931) && !c932) && !c933) && !c934) && !c935) && !c936) && !c937) && !c938) && !c939) && !c940) && !c941) && !c942) && c943); */
          /* c1133 <= ((((((((((((((((((((((((((((!c916 && !c917) && !c918) && !c919) && !c920) && !c921) && !c922) && !c923) && !c924) && !c925) && !c926) && !c927) && !c928) && !c929) && !c930) && !c931) && !c932) && !c933) && !c934) && !c935) && !c936) && !c937) && !c938) && !c939) && !c940) && !c941) && !c942) && !c943) && c944); */
          /* c1134 <= (((((((((((((((((((((((((((((!c916 && !c917) && !c918) && !c919) && !c920) && !c921) && !c922) && !c923) && !c924) && !c925) && !c926) && !c927) && !c928) && !c929) && !c930) && !c931) && !c932) && !c933) && !c934) && !c935) && !c936) && !c937) && !c938) && !c939) && !c940) && !c941) && !c942) && !c943) && !c944) && c945); */
          /* c1135 <= ((((((((((((((((((((((((((((((!c916 && !c917) && !c918) && !c919) && !c920) && !c921) && !c922) && !c923) && !c924) && !c925) && !c926) && !c927) && !c928) && !c929) && !c930) && !c931) && !c932) && !c933) && !c934) && !c935) && !c936) && !c937) && !c938) && !c939) && !c940) && !c941) && !c942) && !c943) && !c944) && !c945) && c946); */
          /* c1136 <= ((((((((((((((((((((((((((((((!c916 && !c917) && !c918) && !c919) && !c920) && !c921) && !c922) && !c923) && !c924) && !c925) && !c926) && !c927) && !c928) && !c929) && !c930) && !c931) && !c932) && !c933) && !c934) && !c935) && !c936) && !c937) && !c938) && !c939) && !c940) && !c941) && !c942) && !c943) && !c944) && !c945) && !c946); */
          if (c916) begin
            a6 <= (c2157 && c916) ? a6 : c2159 ? a6 : c2160 ? a6 : c2161 ? a6 : c2162 ? a6 : c2163 ? a6 : c2164 ? a6 : c2246 ? a6 : c2247 ? a6 : c2166 ? a6 : c2167 ? a6 : c2168 ? stack0_top2 : c2169 ? stack0_top2 : c2170 ? stack0_top2 : c2171 ? stack0_top2 : c2172 ? a6 : c2173 ? a6 : c2174 ? a6 : c2175 ? a6 : c2176 ? a6 : (c2286 || c2284) ? a6 : c2178 ? a6 : c2179 ? a6 : c2180 ? a6 : c2181 ? a6 : c2182 ? a6 : c2212 ? a6 : (c2183 && !c964) ? a6 : c2184 ? a6 : c2185 ? a6 : c2186 ? a6 : c2187 ? a6 : (c2361 || c2360) ? a6 : (c2188 && !c967) ? a6 : (c2157 && c1136) ? a6 : c2158 ? a6 : 'bz;
            /* address0_pos8 <= (c2157 && c916) ? address0_pos2 : c2159 ? address0_pos2 : c2160 ? address0_pos2 : c2161 ? address0_pos2 : c2162 ? address0_pos2 : c2163 ? address0_pos3 : c2164 ? address0_pos4 : c2246 ? address0_pos2 : c2247 ? address0_pos2 : c2166 ? address0_pos2 : c2167 ? address0_pos5 : c2168 ? address0_pos2 : c2169 ? address0_pos2 : c2170 ? address0_pos2 : c2171 ? address0_pos2 : c2172 ? address0_pos2 : c2173 ? address0_pos2 : c2174 ? address0_pos2 : c2175 ? address0_pos2 : c2176 ? address0_pos2 : (c2286 || c2284) ? address0_pos2 : c2178 ? address0_pos2 : c2179 ? address0_pos2 : c2180 ? address0_pos2 : c2181 ? address0_pos2 : c2182 ? address0_pos2 : c2212 ? address0_pos6 : (c2183 && !c964) ? address0_pos2 : c2184 ? address0_pos2 : c2185 ? address0_pos2 : c2186 ? address0_pos2 : c2187 ? address0_pos2 : (c2361 || c2360) ? address0_pos2 : (c2188 && !c967) ? address0_pos2 : (c2157 && c1136) ? address0_pos2 : c2158 ? address0_pos7 : 'bz; */
            /* address0_second8 <= (c2157 && c916) ? address0_second2 : c2159 ? address0_second2 : c2160 ? address0_second2 : c2161 ? address0_second2 : c2162 ? address0_second2 : c2163 ? address0_top2 : c2164 ? address0_second4 : c2246 ? address0_second2 : c2247 ? address0_second2 : c2166 ? address0_second2 : c2167 ? address0_second5 : c2168 ? address0_second2 : c2169 ? address0_second2 : c2170 ? address0_second2 : c2171 ? address0_second2 : c2172 ? address0_second2 : c2173 ? address0_second2 : c2174 ? address0_second2 : c2175 ? address0_second2 : c2176 ? address0_second2 : (c2286 || c2284) ? address0_second2 : c2178 ? address0_second2 : c2179 ? address0_second2 : c2180 ? address0_second2 : c2181 ? address0_second2 : c2182 ? address0_second2 : c2212 ? address0_second6 : (c2183 && !c964) ? address0_second2 : c2184 ? address0_second2 : c2185 ? address0_second2 : c2186 ? address0_second2 : c2187 ? address0_second2 : (c2361 || c2360) ? address0_second2 : (c2188 && !c967) ? address0_second2 : (c2157 && c1136) ? address0_second2 : c2158 ? address0_top2 : 'bz; */
            /* address0_top8 <= (c2157 && c916) ? address0_top2 : c2159 ? address0_top2 : c2160 ? address0_top2 : c2161 ? address0_top2 : c2162 ? address0_top2 : c2163 ? stack0_top2 : c2164 ? address0_second2 : c2246 ? address0_top2 : c2247 ? address0_top2 : c2166 ? address0_top2 : c2167 ? address0_second2 : c2168 ? address0_top2 : c2169 ? address0_top2 : c2170 ? address0_top2 : c2171 ? address0_top2 : c2172 ? address0_top2 : c2173 ? address0_top2 : c2174 ? address0_top2 : c2175 ? address0_top2 : c2176 ? address0_top2 : (c2286 || c2284) ? address0_top2 : c2178 ? address0_top2 : c2179 ? address0_top2 : c2180 ? address0_top2 : c2181 ? address0_top2 : c2182 ? address0_top2 : c2212 ? address0_second2 : (c2183 && !c964) ? address0_top2 : c2184 ? address0_top2 : c2185 ? address0_top2 : c2186 ? address0_top2 : c2187 ? address0_top2 : (c2361 || c2360) ? address0_top2 : (c2188 && !c967) ? address0_top2 : (c2157 && c1136) ? address0_top2 : c2158 ? ip2 : 'bz; */
            b6 <= (c2157 && c916) ? b6 : c2159 ? b6 : c2160 ? b6 : c2161 ? b6 : c2162 ? b6 : c2163 ? b6 : c2164 ? b6 : c2246 ? b6 : c2247 ? b6 : c2166 ? b6 : c2167 ? b6 : c2168 ? stack0_second2 : c2169 ? stack0_second2 : c2170 ? stack0_second2 : c2171 ? stack0_second2 : c2172 ? b6 : c2173 ? b6 : c2174 ? b6 : c2175 ? b6 : c2176 ? b6 : (c2286 || c2284) ? b6 : c2178 ? b6 : c2179 ? b6 : c2180 ? b6 : c2181 ? b6 : c2182 ? b6 : c2212 ? b6 : (c2183 && !c964) ? b6 : c2184 ? b6 : c2185 ? b6 : c2186 ? b6 : c2187 ? b6 : (c2361 || c2360) ? b6 : (c2188 && !c967) ? b6 : (c2157 && c1136) ? b6 : c2158 ? b6 : 'bz;
            /* ip21 <= (c2157 && c916) ? ip2 : c2159 ? ip3 : c2160 ? ip2 : c2161 ? ip2 : c2162 ? ip2 : c2163 ? ip2 : c2164 ? ip2 : c2246 ? ip5 : c2247 ? ip6 : c2166 ? ip8 : c2167 ? address0_top2 : c2168 ? t2660 : c2169 ? t2670 : c2170 ? t2680 : c2171 ? t2690 : c2172 ? ip2 : c2173 ? ip2 : c2174 ? ip2 : c2175 ? ip2 : c2176 ? ip2 : (c2286 || c2284) ? ip2 : c2178 ? ip2 : c2179 ? ip2 : c2180 ? ip2 : c2181 ? ip2 : c2182 ? ip2 : c2212 ? address0_top2 : (c2183 && !c964) ? ip2 : c2184 ? ip2 : c2185 ? ip2 : c2186 ? ip2 : c2187 ? ip2 : (c2361 || c2360) ? ip_inl514 : (c2188 && !c967) ? ip2 : (c2157 && c1136) ? ip2 : c2158 ? ip20 : 'bz; */
            /* stack0_pos35 <= (c2157 && c916) ? stack0_pos2 : c2159 ? stack0_pos3 : c2160 ? stack0_pos4 : c2161 ? stack0_pos5 : c2162 ? stack0_pos2 : c2163 ? stack0_pos6 : c2164 ? stack0_pos7 : c2246 ? stack0_pos2 : c2247 ? stack0_pos8 : c2166 ? stack0_pos2 : c2167 ? stack0_pos2 : c2168 ? stack0_pos10 : c2169 ? stack0_pos12 : c2170 ? stack0_pos14 : c2171 ? stack0_pos16 : c2172 ? stack0_pos2 : c2173 ? stack0_pos18 : c2174 ? stack0_pos19 : c2175 ? stack0_pos20 : c2176 ? stack0_pos21 : (c2286 || c2284) ? stack0_pos2 : c2178 ? stack0_pos22 : c2179 ? stack0_pos23 : c2180 ? stack0_pos24 : c2181 ? stack0_pos25 : c2182 ? stack0_pos26 : c2212 ? stack0_pos27 : (c2183 && !c964) ? stack0_pos2 : c2184 ? stack0_pos2 : c2185 ? stack0_pos2 : c2186 ? stack0_pos2 : c2187 ? stack0_pos29 : (c2361 || c2360) ? stack0_pos34 : (c2188 && !c967) ? stack0_pos2 : (c2157 && c1136) ? stack0_pos2 : c2158 ? stack0_pos2 : 'bz; */
            /* stack0_second37 <= (c2157 && c916) ? stack0_second2 : c2159 ? stack0_top2 : c2160 ? stack0_top2 : c2161 ? stack0_second5 : c2162 ? stack0_top2 : c2163 ? stack0_second7 : c2164 ? stack0_top2 : c2246 ? stack0_second2 : c2247 ? stack0_second9 : c2166 ? stack0_second2 : c2167 ? stack0_second2 : c2168 ? stack0_second11 : c2169 ? stack0_second13 : c2170 ? stack0_second15 : c2171 ? stack0_second17 : c2172 ? stack0_second2 : c2173 ? stack0_second19 : c2174 ? stack0_second20 : c2175 ? stack0_second21 : c2176 ? stack0_second22 : (c2286 || c2284) ? stack0_second23 : c2178 ? stack0_second24 : c2179 ? stack0_second25 : c2180 ? stack0_second26 : c2181 ? stack0_second27 : c2182 ? stack0_second28 : c2212 ? stack0_second29 : (c2183 && !c964) ? stack0_second2 : c2184 ? stack0_second2 : c2185 ? stack0_second2 : c2186 ? stack0_second2 : c2187 ? stack0_second31 : (c2361 || c2360) ? stack0_second36 : (c2188 && !c967) ? stack0_second2 : (c2157 && c1136) ? stack0_second2 : c2158 ? stack0_second2 : 'bz; */
            /* stack0_top50 <= (c2157 && c916) ? stack0_top2 : c2159 ? t947 : c2160 ? stack0_top2 : c2161 ? stack0_second2 : c2162 ? stack0_second2 : c2163 ? stack0_second2 : c2164 ? address0_top2 : c2246 ? stack0_top9 : c2247 ? stack0_second2 : c2166 ? stack0_top2 : c2167 ? stack0_top2 : c2168 ? stack0_second10 : c2169 ? stack0_second12 : c2170 ? stack0_second14 : c2171 ? stack0_second16 : c2172 ? stack0_top19 : c2173 ? stack0_second18 : c2174 ? stack0_top23 : c2175 ? stack0_top25 : c2176 ? stack0_top27 : (c2286 || c2284) ? stack0_top28 : c2178 ? stack0_top30 : c2179 ? stack0_top32 : c2180 ? stack0_top34 : c2181 ? stack0_top36 : c2182 ? stack0_top38 : c2212 ? stack0_second2 : (c2183 && !c964) ? stack0_top2 : c2184 ? stack0_top40 : c2185 ? stack0_top41 : c2186 ? stack0_top42 : c2187 ? stack0_second30 : (c2361 || c2360) ? stack0_top49 : (c2188 && !c967) ? stack0_top2 : (c2157 && c1136) ? stack0_top2 : c2158 ? stack0_top2 : 'bz; */
            t11 <= (c2157 && c916) ? t11 : c2159 ? t11 : c2160 ? t11 : c2161 ? t11 : c2162 ? t11 : c2163 ? t11 : c2164 ? t11 : c2246 ? t11 : c2247 ? t11 : c2166 ? t11 : c2167 ? t11 : c2168 ? t11 : c2169 ? t11 : c2170 ? t11 : c2171 ? t11 : c2172 ? t11 : c2173 ? t11 : c2174 ? stack0_top2 : c2175 ? stack0_top2 : c2176 ? stack0_top2 : (c2286 || c2284) ? t11 : c2178 ? stack0_top2 : c2179 ? stack0_top2 : c2180 ? stack0_top2 : c2181 ? stack0_top2 : c2182 ? stack0_top2 : c2212 ? t11 : (c2183 && !c964) ? t11 : c2184 ? t11 : c2185 ? t11 : c2186 ? stack0_top2 : c2187 ? t11 : (c2361 || c2360) ? t11 : (c2188 && !c967) ? t11 : (c2157 && c1136) ? t11 : c2158 ? t11 : 'bz;
            /* ip22 <= (ip21 + 1); */
            address0_pos2 <= address0_pos8;
            address0_second2 <= address0_second8;
            stack0_pos2 <= stack0_pos35;
            stack0_second2 <= stack0_second37;
            address0_top2 <= address0_top8;
            ip2 <= ip22;
            stack0_top2 <= stack0_top50;
            retro_main_state <= retro_main_L1_b198_S1;
          end else if (c1106) begin
            _stack_addr <= t843_inl3;
            _stack_we <= 1;
            _stack_req <= 1;
            _stack_d <= stack0_second2;
            memory_addr <= ip3;
            memory_we <= 0;
            memory_req <= 1;
            /* ip3 <= (ip2 + 1); */
            /* t843_inl3 <= (stack0_pos2 - 2); */
            /* stack0_pos3 <= (stack0_pos2 + 1); */
            /* c2858 <= (c2856 && c1106); */
            /* c2159 <= (c2157 && c1106); */
            retro_main_state <= retro_main_L1_ifthen11_S1;
          end else if (c1107) begin
            _stack_addr <= t843_inl4;
            _stack_we <= 1;
            _stack_req <= 1;
            _stack_d <= stack0_second2;
            /* t843_inl4 <= (stack0_pos2 - 2); */
            /* stack0_pos4 <= (stack0_pos2 + 1); */
            /* c2859 <= (c2856 && c1107); */
            /* c2160 <= (c2157 && c1107); */
            retro_main_state <= retro_main_L1_ifthen15_S1;
          end else if (c1108) begin
            _stack_addr <= t846_inl8;
            _stack_we <= 0;
            _stack_req <= 1;
            /* stack0_pos5 <= (stack0_pos2 - 1); */
            /* t846_inl8 <= (stack0_pos5 - 2); */
            /* c2860 <= (c2856 && c1108); */
            /* c2161 <= (c2157 && c1108); */
            retro_main_state <= retro_main_L1_ifthen19_S1;
          end else if (c1109) begin
            /* c2861 <= (c2856 && c1109); */
            /* c2162 <= (c2157 && c1109); */
            retro_main_state <= retro_main_L1_b198_S0;
          end else if (c1110) begin
            _stack_addr <= t846_inl9;
            _stack_we <= 0;
            _stack_req <= 1;
            _address_addr <= t843_inl5;
            _address_we <= 1;
            _address_req <= 1;
            _address_d <= address0_second2;
            /* stack0_pos6 <= (stack0_pos2 - 1); */
            /* t843_inl5 <= (address0_pos2 - 2); */
            /* address0_pos3 <= (address0_pos2 + 1); */
            /* t846_inl9 <= (stack0_pos6 - 2); */
            /* c2862 <= (c2856 && c1110); */
            /* c2163 <= (c2157 && c1110); */
            retro_main_state <= retro_main_L1_ifthen27_S1;
          end else if (c1111) begin
            _address_addr <= t846_inl10;
            _address_we <= 0;
            _address_req <= 1;
            _stack_addr <= t843_inl6;
            _stack_we <= 1;
            _stack_req <= 1;
            _stack_d <= stack0_second2;
            /* address0_pos4 <= (address0_pos2 - 1); */
            /* t843_inl6 <= (stack0_pos2 - 2); */
            /* stack0_pos7 <= (stack0_pos2 + 1); */
            /* t846_inl10 <= (address0_pos4 - 2); */
            /* c2863 <= (c2856 && c1111); */
            /* c2164 <= (c2157 && c1111); */
            retro_main_state <= retro_main_L1_ifthen31_S1;
          end else if (c1112) begin
            /* stack0_top9 <= (stack0_top2 - 1); */
            /* c950 <= (stack0_top9 != 0); */
            /* c951 <= (stack0_top9 > -1); */
            /* c952 <= (c950 && c951); */
            /* c2864 <= (c2856 && c1112); */
            /* c2165 <= (c2157 && c1112); */
            if (c952) begin
              memory_addr <= ip4;
              memory_we <= 0;
              memory_req <= 1;
              /* ip4 <= (ip2 + 1); */
              /* c2888 <= (c2864 && c952); */
              /* c2246 <= (c2165 && c952); */
              retro_main_state <= retro_main_L1_ifthen38_S1;
            end else begin
              _stack_addr <= t846_inl11;
              _stack_we <= 0;
              _stack_req <= 1;
              /* ip6 <= (ip2 + 1); */
              /* stack0_pos8 <= (stack0_pos2 - 1); */
              /* t846_inl11 <= (stack0_pos8 - 2); */
              /* c2889 <= (c2864 && !c952); */
              /* c2247 <= (c2165 && !c952); */
              retro_main_state <= retro_main_L1_ifelse41_S1;
            end
          end else if (c1113) begin
            memory_addr <= ip7;
            memory_we <= 0;
            memory_req <= 1;
            /* ip7 <= (ip2 + 1); */
            /* c2865 <= (c2856 && c1113); */
            /* c2166 <= (c2157 && c1113); */
            retro_main_state <= retro_main_L1_ifthen44_S1;
          end else if (c1114) begin
            _address_addr <= t846_inl12;
            _address_we <= 0;
            _address_req <= 1;
            /* address0_pos5 <= (address0_pos2 - 1); */
            /* t846_inl12 <= (address0_pos5 - 2); */
            /* c2866 <= (c2856 && c1114); */
            /* c2167 <= (c2157 && c1114); */
            retro_main_state <= retro_main_L1_ifthen48_S1;
          end else if (c1115) begin
            _stack_addr <= t846_inl13;
            _stack_we <= 0;
            _stack_req <= 1;
            /* ip10 <= (ip2 + 1); */
            /* stack0_pos9 <= (stack0_pos2 - 1); */
            /* c955 <= (stack0_second2 > stack0_top2); */
            /* t846_inl13 <= (stack0_pos9 - 2); */
            /* stack0_pos10 <= (stack0_pos9 - 1); */
            /* t846_inl14 <= (stack0_pos10 - 2); */
            /* c2867 <= (c2856 && c1115); */
            /* c2168 <= (c2157 && c1115); */
            /* c2277 <= (c2168 && c955); */
            retro_main_state <= retro_main_L1_ifthen52_S1;
          end else if (c1116) begin
            _stack_addr <= t846_inl15;
            _stack_we <= 0;
            _stack_req <= 1;
            /* ip12 <= (ip2 + 1); */
            /* stack0_pos11 <= (stack0_pos2 - 1); */
            /* c957 <= (stack0_second2 < stack0_top2); */
            /* t846_inl15 <= (stack0_pos11 - 2); */
            /* stack0_pos12 <= (stack0_pos11 - 1); */
            /* t846_inl16 <= (stack0_pos12 - 2); */
            /* c2868 <= (c2856 && c1116); */
            /* c2169 <= (c2157 && c1116); */
            /* c2278 <= (c2169 && c957); */
            retro_main_state <= retro_main_L1_ifthen61_S1;
          end else if (c1117) begin
            _stack_addr <= t846_inl17;
            _stack_we <= 0;
            _stack_req <= 1;
            /* ip14 <= (ip2 + 1); */
            /* stack0_pos13 <= (stack0_pos2 - 1); */
            /* c959 <= (stack0_second2 != stack0_top2); */
            /* t846_inl17 <= (stack0_pos13 - 2); */
            /* stack0_pos14 <= (stack0_pos13 - 1); */
            /* t846_inl18 <= (stack0_pos14 - 2); */
            /* c2869 <= (c2856 && c1117); */
            /* c2170 <= (c2157 && c1117); */
            /* c2279 <= (c2170 && c959); */
            retro_main_state <= retro_main_L1_ifthen70_S1;
          end else if (c1118) begin
            _stack_addr <= t846_inl19;
            _stack_we <= 0;
            _stack_req <= 1;
            /* ip16 <= (ip2 + 1); */
            /* stack0_pos15 <= (stack0_pos2 - 1); */
            /* c961 <= (stack0_second2 == stack0_top2); */
            /* t846_inl19 <= (stack0_pos15 - 2); */
            /* stack0_pos16 <= (stack0_pos15 - 1); */
            /* t846_inl20 <= (stack0_pos16 - 2); */
            /* c2870 <= (c2856 && c1118); */
            /* c2171 <= (c2157 && c1118); */
            /* c2280 <= (c2171 && c961); */
            retro_main_state <= retro_main_L1_ifthen79_S1;
          end else if (c1119) begin
            memory_addr <= stack0_top2;
            memory_we <= 0;
            memory_req <= 1;
            /* c2871 <= (c2856 && c1119); */
            /* c2172 <= (c2157 && c1119); */
            retro_main_state <= retro_main_L1_ifthen88_S1;
          end else if (c1120) begin
            _stack_addr <= t846_inl21;
            _stack_we <= 0;
            _stack_req <= 1;
            memory_addr <= stack0_top2;
            memory_we <= 1;
            memory_req <= 1;
            memory_d <= stack0_second2;
            /* stack0_pos17 <= (stack0_pos2 - 1); */
            /* t846_inl21 <= (stack0_pos17 - 2); */
            /* stack0_pos18 <= (stack0_pos17 - 1); */
            /* t846_inl22 <= (stack0_pos18 - 2); */
            /* c2872 <= (c2856 && c1120); */
            /* c2173 <= (c2157 && c1120); */
            retro_main_state <= retro_main_L1_ifthen92_S1;
          end else if (c1121) begin
            _stack_addr <= t846_inl23;
            _stack_we <= 0;
            _stack_req <= 1;
            /* stack0_pos19 <= (stack0_pos2 - 1); */
            /* stack0_top23 <= (stack0_second2 + stack0_top2); */
            /* t846_inl23 <= (stack0_pos19 - 2); */
            /* c2873 <= (c2856 && c1121); */
            /* c2174 <= (c2157 && c1121); */
            retro_main_state <= retro_main_L1_ifthen96_S1;
          end else if (c1122) begin
            _stack_addr <= t846_inl24;
            _stack_we <= 0;
            _stack_req <= 1;
            /* stack0_pos20 <= (stack0_pos2 - 1); */
            /* stack0_top25 <= (stack0_second2 - stack0_top2); */
            /* t846_inl24 <= (stack0_pos20 - 2); */
            /* c2874 <= (c2856 && c1122); */
            /* c2175 <= (c2157 && c1122); */
            retro_main_state <= retro_main_L1_ifthen100_S1;
          end else if (c1123) begin
            _stack_addr <= t846_inl25;
            _stack_we <= 0;
            _stack_req <= 1;
            /* stack0_pos21 <= (stack0_pos2 - 1); */
            /* stack0_top27 <= (stack0_second2 * stack0_top2); */
            /* t846_inl25 <= (stack0_pos21 - 2); */
            /* c2875 <= (c2856 && c1123); */
            /* c2176 <= (c2157 && c1123); */
            retro_main_state <= retro_main_L1_ifthen104_S1;
          end else if (c1124) begin
            /* t969_inl49 <= (stack0_second2 & 2147483648); */
            /* t971_inl49 <= (stack0_top2 & 2147483648); */
            /* abs_a_inl492 <= (stack0_second2 & 2147483647); */
            /* abs_b_inl492 <= (stack0_top2 & 2147483647); */
            i_inl1_inl493 <= 0;
            n_inl1_inl493 <= 0;
            test_bit_inl1_inl493 <= 1073741824;
            /* t970_inl49 <= t969_inl49 ? 1 : 0; */
            /* t972_inl49 <= t971_inl49 ? 1 : 0; */
            /* x_inl1_inl49 <= abs_a_inl492; */
            /* c2876 <= (c2856 && c1124); */
            /* c2177 <= (c2157 && c1124); */
            retro_main_state <= retro_main_L20_fortest393_S0;
          end else if (c1125) begin
            _stack_addr <= t846_inl26;
            _stack_we <= 0;
            _stack_req <= 1;
            /* stack0_pos22 <= (stack0_pos2 - 1); */
            /* stack0_top30 <= (stack0_second2 & stack0_top2); */
            /* t846_inl26 <= (stack0_pos22 - 2); */
            /* c2877 <= (c2856 && c1125); */
            /* c2178 <= (c2157 && c1125); */
            retro_main_state <= retro_main_L1_ifthen112_S1;
          end else if (c1126) begin
            _stack_addr <= t846_inl27;
            _stack_we <= 0;
            _stack_req <= 1;
            /* stack0_pos23 <= (stack0_pos2 - 1); */
            /* stack0_top32 <= (stack0_second2 | stack0_top2); */
            /* t846_inl27 <= (stack0_pos23 - 2); */
            /* c2878 <= (c2856 && c1126); */
            /* c2179 <= (c2157 && c1126); */
            retro_main_state <= retro_main_L1_ifthen116_S1;
          end else if (c1127) begin
            _stack_addr <= t846_inl28;
            _stack_we <= 0;
            _stack_req <= 1;
            /* stack0_pos24 <= (stack0_pos2 - 1); */
            /* stack0_top34 <= (stack0_second2 ^ stack0_top2); */
            /* t846_inl28 <= (stack0_pos24 - 2); */
            /* c2879 <= (c2856 && c1127); */
            /* c2180 <= (c2157 && c1127); */
            retro_main_state <= retro_main_L1_ifthen120_S1;
          end else if (c1128) begin
            _stack_addr <= t846_inl29;
            _stack_we <= 0;
            _stack_req <= 1;
            /* stack0_pos25 <= (stack0_pos2 - 1); */
            /* stack0_top36 <= (stack0_second2 << stack0_top2); */
            /* t846_inl29 <= (stack0_pos25 - 2); */
            /* c2880 <= (c2856 && c1128); */
            /* c2181 <= (c2157 && c1128); */
            retro_main_state <= retro_main_L1_ifthen124_S1;
          end else if (c1129) begin
            _stack_addr <= t846_inl30;
            _stack_we <= 0;
            _stack_req <= 1;
            /* stack0_pos26 <= (stack0_pos2 - 1); */
            /* stack0_top38 <= (stack0_second2 >>> stack0_top2); */
            /* t846_inl30 <= (stack0_pos26 - 2); */
            /* c2881 <= (c2856 && c1129); */
            /* c2182 <= (c2157 && c1129); */
            retro_main_state <= retro_main_L1_ifthen128_S1;
          end else if (c1130) begin
            /* c964 <= (stack0_top2 == 0); */
            /* c2882 <= (c2856 && c1130); */
            /* c2183 <= (c2157 && c1130); */
            if (c964) begin
              _address_addr <= t846_inl32;
              _address_we <= 0;
              _address_req <= 1;
              _stack_addr <= t846_inl31;
              _stack_we <= 0;
              _stack_req <= 1;
              /* stack0_pos27 <= (stack0_pos2 - 1); */
              /* address0_pos6 <= (address0_pos2 - 1); */
              /* t846_inl31 <= (stack0_pos27 - 2); */
              /* t846_inl32 <= (address0_pos6 - 2); */
              /* c2894 <= (c2882 && c964); */
              /* c2212 <= (c2183 && c964); */
              retro_main_state <= retro_main_L1_ifthen135_S1;
            end else begin
              a6 <= (c2157 && c916) ? a6 : c2159 ? a6 : c2160 ? a6 : c2161 ? a6 : c2162 ? a6 : c2163 ? a6 : c2164 ? a6 : c2246 ? a6 : c2247 ? a6 : c2166 ? a6 : c2167 ? a6 : c2168 ? stack0_top2 : c2169 ? stack0_top2 : c2170 ? stack0_top2 : c2171 ? stack0_top2 : c2172 ? a6 : c2173 ? a6 : c2174 ? a6 : c2175 ? a6 : c2176 ? a6 : (c2286 || c2284) ? a6 : c2178 ? a6 : c2179 ? a6 : c2180 ? a6 : c2181 ? a6 : c2182 ? a6 : c2212 ? a6 : (c2183 && !c964) ? a6 : c2184 ? a6 : c2185 ? a6 : c2186 ? a6 : c2187 ? a6 : (c2361 || c2360) ? a6 : (c2188 && !c967) ? a6 : (c2157 && c1136) ? a6 : c2158 ? a6 : 'bz;
              /* address0_pos8 <= (c2157 && c916) ? address0_pos2 : c2159 ? address0_pos2 : c2160 ? address0_pos2 : c2161 ? address0_pos2 : c2162 ? address0_pos2 : c2163 ? address0_pos3 : c2164 ? address0_pos4 : c2246 ? address0_pos2 : c2247 ? address0_pos2 : c2166 ? address0_pos2 : c2167 ? address0_pos5 : c2168 ? address0_pos2 : c2169 ? address0_pos2 : c2170 ? address0_pos2 : c2171 ? address0_pos2 : c2172 ? address0_pos2 : c2173 ? address0_pos2 : c2174 ? address0_pos2 : c2175 ? address0_pos2 : c2176 ? address0_pos2 : (c2286 || c2284) ? address0_pos2 : c2178 ? address0_pos2 : c2179 ? address0_pos2 : c2180 ? address0_pos2 : c2181 ? address0_pos2 : c2182 ? address0_pos2 : c2212 ? address0_pos6 : (c2183 && !c964) ? address0_pos2 : c2184 ? address0_pos2 : c2185 ? address0_pos2 : c2186 ? address0_pos2 : c2187 ? address0_pos2 : (c2361 || c2360) ? address0_pos2 : (c2188 && !c967) ? address0_pos2 : (c2157 && c1136) ? address0_pos2 : c2158 ? address0_pos7 : 'bz; */
              /* address0_second8 <= (c2157 && c916) ? address0_second2 : c2159 ? address0_second2 : c2160 ? address0_second2 : c2161 ? address0_second2 : c2162 ? address0_second2 : c2163 ? address0_top2 : c2164 ? address0_second4 : c2246 ? address0_second2 : c2247 ? address0_second2 : c2166 ? address0_second2 : c2167 ? address0_second5 : c2168 ? address0_second2 : c2169 ? address0_second2 : c2170 ? address0_second2 : c2171 ? address0_second2 : c2172 ? address0_second2 : c2173 ? address0_second2 : c2174 ? address0_second2 : c2175 ? address0_second2 : c2176 ? address0_second2 : (c2286 || c2284) ? address0_second2 : c2178 ? address0_second2 : c2179 ? address0_second2 : c2180 ? address0_second2 : c2181 ? address0_second2 : c2182 ? address0_second2 : c2212 ? address0_second6 : (c2183 && !c964) ? address0_second2 : c2184 ? address0_second2 : c2185 ? address0_second2 : c2186 ? address0_second2 : c2187 ? address0_second2 : (c2361 || c2360) ? address0_second2 : (c2188 && !c967) ? address0_second2 : (c2157 && c1136) ? address0_second2 : c2158 ? address0_top2 : 'bz; */
              /* address0_top8 <= (c2157 && c916) ? address0_top2 : c2159 ? address0_top2 : c2160 ? address0_top2 : c2161 ? address0_top2 : c2162 ? address0_top2 : c2163 ? stack0_top2 : c2164 ? address0_second2 : c2246 ? address0_top2 : c2247 ? address0_top2 : c2166 ? address0_top2 : c2167 ? address0_second2 : c2168 ? address0_top2 : c2169 ? address0_top2 : c2170 ? address0_top2 : c2171 ? address0_top2 : c2172 ? address0_top2 : c2173 ? address0_top2 : c2174 ? address0_top2 : c2175 ? address0_top2 : c2176 ? address0_top2 : (c2286 || c2284) ? address0_top2 : c2178 ? address0_top2 : c2179 ? address0_top2 : c2180 ? address0_top2 : c2181 ? address0_top2 : c2182 ? address0_top2 : c2212 ? address0_second2 : (c2183 && !c964) ? address0_top2 : c2184 ? address0_top2 : c2185 ? address0_top2 : c2186 ? address0_top2 : c2187 ? address0_top2 : (c2361 || c2360) ? address0_top2 : (c2188 && !c967) ? address0_top2 : (c2157 && c1136) ? address0_top2 : c2158 ? ip2 : 'bz; */
              b6 <= (c2157 && c916) ? b6 : c2159 ? b6 : c2160 ? b6 : c2161 ? b6 : c2162 ? b6 : c2163 ? b6 : c2164 ? b6 : c2246 ? b6 : c2247 ? b6 : c2166 ? b6 : c2167 ? b6 : c2168 ? stack0_second2 : c2169 ? stack0_second2 : c2170 ? stack0_second2 : c2171 ? stack0_second2 : c2172 ? b6 : c2173 ? b6 : c2174 ? b6 : c2175 ? b6 : c2176 ? b6 : (c2286 || c2284) ? b6 : c2178 ? b6 : c2179 ? b6 : c2180 ? b6 : c2181 ? b6 : c2182 ? b6 : c2212 ? b6 : (c2183 && !c964) ? b6 : c2184 ? b6 : c2185 ? b6 : c2186 ? b6 : c2187 ? b6 : (c2361 || c2360) ? b6 : (c2188 && !c967) ? b6 : (c2157 && c1136) ? b6 : c2158 ? b6 : 'bz;
              /* ip21 <= (c2157 && c916) ? ip2 : c2159 ? ip3 : c2160 ? ip2 : c2161 ? ip2 : c2162 ? ip2 : c2163 ? ip2 : c2164 ? ip2 : c2246 ? ip5 : c2247 ? ip6 : c2166 ? ip8 : c2167 ? address0_top2 : c2168 ? t2660 : c2169 ? t2670 : c2170 ? t2680 : c2171 ? t2690 : c2172 ? ip2 : c2173 ? ip2 : c2174 ? ip2 : c2175 ? ip2 : c2176 ? ip2 : (c2286 || c2284) ? ip2 : c2178 ? ip2 : c2179 ? ip2 : c2180 ? ip2 : c2181 ? ip2 : c2182 ? ip2 : c2212 ? address0_top2 : (c2183 && !c964) ? ip2 : c2184 ? ip2 : c2185 ? ip2 : c2186 ? ip2 : c2187 ? ip2 : (c2361 || c2360) ? ip_inl514 : (c2188 && !c967) ? ip2 : (c2157 && c1136) ? ip2 : c2158 ? ip20 : 'bz; */
              /* stack0_pos35 <= (c2157 && c916) ? stack0_pos2 : c2159 ? stack0_pos3 : c2160 ? stack0_pos4 : c2161 ? stack0_pos5 : c2162 ? stack0_pos2 : c2163 ? stack0_pos6 : c2164 ? stack0_pos7 : c2246 ? stack0_pos2 : c2247 ? stack0_pos8 : c2166 ? stack0_pos2 : c2167 ? stack0_pos2 : c2168 ? stack0_pos10 : c2169 ? stack0_pos12 : c2170 ? stack0_pos14 : c2171 ? stack0_pos16 : c2172 ? stack0_pos2 : c2173 ? stack0_pos18 : c2174 ? stack0_pos19 : c2175 ? stack0_pos20 : c2176 ? stack0_pos21 : (c2286 || c2284) ? stack0_pos2 : c2178 ? stack0_pos22 : c2179 ? stack0_pos23 : c2180 ? stack0_pos24 : c2181 ? stack0_pos25 : c2182 ? stack0_pos26 : c2212 ? stack0_pos27 : (c2183 && !c964) ? stack0_pos2 : c2184 ? stack0_pos2 : c2185 ? stack0_pos2 : c2186 ? stack0_pos2 : c2187 ? stack0_pos29 : (c2361 || c2360) ? stack0_pos34 : (c2188 && !c967) ? stack0_pos2 : (c2157 && c1136) ? stack0_pos2 : c2158 ? stack0_pos2 : 'bz; */
              /* stack0_second37 <= (c2157 && c916) ? stack0_second2 : c2159 ? stack0_top2 : c2160 ? stack0_top2 : c2161 ? stack0_second5 : c2162 ? stack0_top2 : c2163 ? stack0_second7 : c2164 ? stack0_top2 : c2246 ? stack0_second2 : c2247 ? stack0_second9 : c2166 ? stack0_second2 : c2167 ? stack0_second2 : c2168 ? stack0_second11 : c2169 ? stack0_second13 : c2170 ? stack0_second15 : c2171 ? stack0_second17 : c2172 ? stack0_second2 : c2173 ? stack0_second19 : c2174 ? stack0_second20 : c2175 ? stack0_second21 : c2176 ? stack0_second22 : (c2286 || c2284) ? stack0_second23 : c2178 ? stack0_second24 : c2179 ? stack0_second25 : c2180 ? stack0_second26 : c2181 ? stack0_second27 : c2182 ? stack0_second28 : c2212 ? stack0_second29 : (c2183 && !c964) ? stack0_second2 : c2184 ? stack0_second2 : c2185 ? stack0_second2 : c2186 ? stack0_second2 : c2187 ? stack0_second31 : (c2361 || c2360) ? stack0_second36 : (c2188 && !c967) ? stack0_second2 : (c2157 && c1136) ? stack0_second2 : c2158 ? stack0_second2 : 'bz; */
              /* stack0_top50 <= (c2157 && c916) ? stack0_top2 : c2159 ? t947 : c2160 ? stack0_top2 : c2161 ? stack0_second2 : c2162 ? stack0_second2 : c2163 ? stack0_second2 : c2164 ? address0_top2 : c2246 ? stack0_top9 : c2247 ? stack0_second2 : c2166 ? stack0_top2 : c2167 ? stack0_top2 : c2168 ? stack0_second10 : c2169 ? stack0_second12 : c2170 ? stack0_second14 : c2171 ? stack0_second16 : c2172 ? stack0_top19 : c2173 ? stack0_second18 : c2174 ? stack0_top23 : c2175 ? stack0_top25 : c2176 ? stack0_top27 : (c2286 || c2284) ? stack0_top28 : c2178 ? stack0_top30 : c2179 ? stack0_top32 : c2180 ? stack0_top34 : c2181 ? stack0_top36 : c2182 ? stack0_top38 : c2212 ? stack0_second2 : (c2183 && !c964) ? stack0_top2 : c2184 ? stack0_top40 : c2185 ? stack0_top41 : c2186 ? stack0_top42 : c2187 ? stack0_second30 : (c2361 || c2360) ? stack0_top49 : (c2188 && !c967) ? stack0_top2 : (c2157 && c1136) ? stack0_top2 : c2158 ? stack0_top2 : 'bz; */
              t11 <= (c2157 && c916) ? t11 : c2159 ? t11 : c2160 ? t11 : c2161 ? t11 : c2162 ? t11 : c2163 ? t11 : c2164 ? t11 : c2246 ? t11 : c2247 ? t11 : c2166 ? t11 : c2167 ? t11 : c2168 ? t11 : c2169 ? t11 : c2170 ? t11 : c2171 ? t11 : c2172 ? t11 : c2173 ? t11 : c2174 ? stack0_top2 : c2175 ? stack0_top2 : c2176 ? stack0_top2 : (c2286 || c2284) ? t11 : c2178 ? stack0_top2 : c2179 ? stack0_top2 : c2180 ? stack0_top2 : c2181 ? stack0_top2 : c2182 ? stack0_top2 : c2212 ? t11 : (c2183 && !c964) ? t11 : c2184 ? t11 : c2185 ? t11 : c2186 ? stack0_top2 : c2187 ? t11 : (c2361 || c2360) ? t11 : (c2188 && !c967) ? t11 : (c2157 && c1136) ? t11 : c2158 ? t11 : 'bz;
              /* ip22 <= (ip21 + 1); */
              address0_pos2 <= address0_pos8;
              address0_second2 <= address0_second8;
              stack0_pos2 <= stack0_pos35;
              stack0_second2 <= stack0_second37;
              address0_top2 <= address0_top8;
              ip2 <= ip22;
              stack0_top2 <= stack0_top50;
              retro_main_state <= retro_main_L1_b198_S1;
            end
          end else if (c1131) begin
            /* stack0_top40 <= (stack0_top2 + 1); */
            /* c2883 <= (c2856 && c1131); */
            /* c2184 <= (c2157 && c1131); */
            retro_main_state <= retro_main_L1_b198_S0;
          end else if (c1132) begin
            /* stack0_top41 <= (stack0_top2 - 1); */
            /* c2884 <= (c2856 && c1132); */
            /* c2185 <= (c2157 && c1132); */
            retro_main_state <= retro_main_L1_b198_S0;
          end else if (c1133) begin
            stack0_top42 <= array998[stack0_top2];
            array998[stack0_top2] <= 0;
            /* c2885 <= (c2856 && c1133); */
            /* c2186 <= (c2157 && c1133); */
            retro_main_state <= retro_main_L1_b198_S0;
          end else if (c1134) begin
            _stack_addr <= t846_inl33;
            _stack_we <= 0;
            _stack_req <= 1;
            /* stack0_pos28 <= (stack0_pos2 - 1); */
            array998[stack0_top2] <= stack0_second2;
            /* t846_inl33 <= (stack0_pos28 - 2); */
            /* stack0_pos29 <= (stack0_pos28 - 1); */
            /* t846_inl34 <= (stack0_pos29 - 2); */
            /* c2886 <= (c2856 && c1134); */
            /* c2187 <= (c2157 && c1134); */
            retro_main_state <= retro_main_L1_ifthen153_S1;
          end else if (c1135) begin
            t966 <= array998[0];
            /* c2887 <= (c2856 && c1135); */
            /* c2188 <= (c2157 && c1135); */
            retro_main_state <= retro_main_L1_ifthen157_S1;
          end else if (c1136) begin
            a6 <= (c2157 && c916) ? a6 : c2159 ? a6 : c2160 ? a6 : c2161 ? a6 : c2162 ? a6 : c2163 ? a6 : c2164 ? a6 : c2246 ? a6 : c2247 ? a6 : c2166 ? a6 : c2167 ? a6 : c2168 ? stack0_top2 : c2169 ? stack0_top2 : c2170 ? stack0_top2 : c2171 ? stack0_top2 : c2172 ? a6 : c2173 ? a6 : c2174 ? a6 : c2175 ? a6 : c2176 ? a6 : (c2286 || c2284) ? a6 : c2178 ? a6 : c2179 ? a6 : c2180 ? a6 : c2181 ? a6 : c2182 ? a6 : c2212 ? a6 : (c2183 && !c964) ? a6 : c2184 ? a6 : c2185 ? a6 : c2186 ? a6 : c2187 ? a6 : (c2361 || c2360) ? a6 : (c2188 && !c967) ? a6 : (c2157 && c1136) ? a6 : c2158 ? a6 : 'bz;
            /* address0_pos8 <= (c2157 && c916) ? address0_pos2 : c2159 ? address0_pos2 : c2160 ? address0_pos2 : c2161 ? address0_pos2 : c2162 ? address0_pos2 : c2163 ? address0_pos3 : c2164 ? address0_pos4 : c2246 ? address0_pos2 : c2247 ? address0_pos2 : c2166 ? address0_pos2 : c2167 ? address0_pos5 : c2168 ? address0_pos2 : c2169 ? address0_pos2 : c2170 ? address0_pos2 : c2171 ? address0_pos2 : c2172 ? address0_pos2 : c2173 ? address0_pos2 : c2174 ? address0_pos2 : c2175 ? address0_pos2 : c2176 ? address0_pos2 : (c2286 || c2284) ? address0_pos2 : c2178 ? address0_pos2 : c2179 ? address0_pos2 : c2180 ? address0_pos2 : c2181 ? address0_pos2 : c2182 ? address0_pos2 : c2212 ? address0_pos6 : (c2183 && !c964) ? address0_pos2 : c2184 ? address0_pos2 : c2185 ? address0_pos2 : c2186 ? address0_pos2 : c2187 ? address0_pos2 : (c2361 || c2360) ? address0_pos2 : (c2188 && !c967) ? address0_pos2 : (c2157 && c1136) ? address0_pos2 : c2158 ? address0_pos7 : 'bz; */
            /* address0_second8 <= (c2157 && c916) ? address0_second2 : c2159 ? address0_second2 : c2160 ? address0_second2 : c2161 ? address0_second2 : c2162 ? address0_second2 : c2163 ? address0_top2 : c2164 ? address0_second4 : c2246 ? address0_second2 : c2247 ? address0_second2 : c2166 ? address0_second2 : c2167 ? address0_second5 : c2168 ? address0_second2 : c2169 ? address0_second2 : c2170 ? address0_second2 : c2171 ? address0_second2 : c2172 ? address0_second2 : c2173 ? address0_second2 : c2174 ? address0_second2 : c2175 ? address0_second2 : c2176 ? address0_second2 : (c2286 || c2284) ? address0_second2 : c2178 ? address0_second2 : c2179 ? address0_second2 : c2180 ? address0_second2 : c2181 ? address0_second2 : c2182 ? address0_second2 : c2212 ? address0_second6 : (c2183 && !c964) ? address0_second2 : c2184 ? address0_second2 : c2185 ? address0_second2 : c2186 ? address0_second2 : c2187 ? address0_second2 : (c2361 || c2360) ? address0_second2 : (c2188 && !c967) ? address0_second2 : (c2157 && c1136) ? address0_second2 : c2158 ? address0_top2 : 'bz; */
            /* address0_top8 <= (c2157 && c916) ? address0_top2 : c2159 ? address0_top2 : c2160 ? address0_top2 : c2161 ? address0_top2 : c2162 ? address0_top2 : c2163 ? stack0_top2 : c2164 ? address0_second2 : c2246 ? address0_top2 : c2247 ? address0_top2 : c2166 ? address0_top2 : c2167 ? address0_second2 : c2168 ? address0_top2 : c2169 ? address0_top2 : c2170 ? address0_top2 : c2171 ? address0_top2 : c2172 ? address0_top2 : c2173 ? address0_top2 : c2174 ? address0_top2 : c2175 ? address0_top2 : c2176 ? address0_top2 : (c2286 || c2284) ? address0_top2 : c2178 ? address0_top2 : c2179 ? address0_top2 : c2180 ? address0_top2 : c2181 ? address0_top2 : c2182 ? address0_top2 : c2212 ? address0_second2 : (c2183 && !c964) ? address0_top2 : c2184 ? address0_top2 : c2185 ? address0_top2 : c2186 ? address0_top2 : c2187 ? address0_top2 : (c2361 || c2360) ? address0_top2 : (c2188 && !c967) ? address0_top2 : (c2157 && c1136) ? address0_top2 : c2158 ? ip2 : 'bz; */
            b6 <= (c2157 && c916) ? b6 : c2159 ? b6 : c2160 ? b6 : c2161 ? b6 : c2162 ? b6 : c2163 ? b6 : c2164 ? b6 : c2246 ? b6 : c2247 ? b6 : c2166 ? b6 : c2167 ? b6 : c2168 ? stack0_second2 : c2169 ? stack0_second2 : c2170 ? stack0_second2 : c2171 ? stack0_second2 : c2172 ? b6 : c2173 ? b6 : c2174 ? b6 : c2175 ? b6 : c2176 ? b6 : (c2286 || c2284) ? b6 : c2178 ? b6 : c2179 ? b6 : c2180 ? b6 : c2181 ? b6 : c2182 ? b6 : c2212 ? b6 : (c2183 && !c964) ? b6 : c2184 ? b6 : c2185 ? b6 : c2186 ? b6 : c2187 ? b6 : (c2361 || c2360) ? b6 : (c2188 && !c967) ? b6 : (c2157 && c1136) ? b6 : c2158 ? b6 : 'bz;
            /* ip21 <= (c2157 && c916) ? ip2 : c2159 ? ip3 : c2160 ? ip2 : c2161 ? ip2 : c2162 ? ip2 : c2163 ? ip2 : c2164 ? ip2 : c2246 ? ip5 : c2247 ? ip6 : c2166 ? ip8 : c2167 ? address0_top2 : c2168 ? t2660 : c2169 ? t2670 : c2170 ? t2680 : c2171 ? t2690 : c2172 ? ip2 : c2173 ? ip2 : c2174 ? ip2 : c2175 ? ip2 : c2176 ? ip2 : (c2286 || c2284) ? ip2 : c2178 ? ip2 : c2179 ? ip2 : c2180 ? ip2 : c2181 ? ip2 : c2182 ? ip2 : c2212 ? address0_top2 : (c2183 && !c964) ? ip2 : c2184 ? ip2 : c2185 ? ip2 : c2186 ? ip2 : c2187 ? ip2 : (c2361 || c2360) ? ip_inl514 : (c2188 && !c967) ? ip2 : (c2157 && c1136) ? ip2 : c2158 ? ip20 : 'bz; */
            /* stack0_pos35 <= (c2157 && c916) ? stack0_pos2 : c2159 ? stack0_pos3 : c2160 ? stack0_pos4 : c2161 ? stack0_pos5 : c2162 ? stack0_pos2 : c2163 ? stack0_pos6 : c2164 ? stack0_pos7 : c2246 ? stack0_pos2 : c2247 ? stack0_pos8 : c2166 ? stack0_pos2 : c2167 ? stack0_pos2 : c2168 ? stack0_pos10 : c2169 ? stack0_pos12 : c2170 ? stack0_pos14 : c2171 ? stack0_pos16 : c2172 ? stack0_pos2 : c2173 ? stack0_pos18 : c2174 ? stack0_pos19 : c2175 ? stack0_pos20 : c2176 ? stack0_pos21 : (c2286 || c2284) ? stack0_pos2 : c2178 ? stack0_pos22 : c2179 ? stack0_pos23 : c2180 ? stack0_pos24 : c2181 ? stack0_pos25 : c2182 ? stack0_pos26 : c2212 ? stack0_pos27 : (c2183 && !c964) ? stack0_pos2 : c2184 ? stack0_pos2 : c2185 ? stack0_pos2 : c2186 ? stack0_pos2 : c2187 ? stack0_pos29 : (c2361 || c2360) ? stack0_pos34 : (c2188 && !c967) ? stack0_pos2 : (c2157 && c1136) ? stack0_pos2 : c2158 ? stack0_pos2 : 'bz; */
            /* stack0_second37 <= (c2157 && c916) ? stack0_second2 : c2159 ? stack0_top2 : c2160 ? stack0_top2 : c2161 ? stack0_second5 : c2162 ? stack0_top2 : c2163 ? stack0_second7 : c2164 ? stack0_top2 : c2246 ? stack0_second2 : c2247 ? stack0_second9 : c2166 ? stack0_second2 : c2167 ? stack0_second2 : c2168 ? stack0_second11 : c2169 ? stack0_second13 : c2170 ? stack0_second15 : c2171 ? stack0_second17 : c2172 ? stack0_second2 : c2173 ? stack0_second19 : c2174 ? stack0_second20 : c2175 ? stack0_second21 : c2176 ? stack0_second22 : (c2286 || c2284) ? stack0_second23 : c2178 ? stack0_second24 : c2179 ? stack0_second25 : c2180 ? stack0_second26 : c2181 ? stack0_second27 : c2182 ? stack0_second28 : c2212 ? stack0_second29 : (c2183 && !c964) ? stack0_second2 : c2184 ? stack0_second2 : c2185 ? stack0_second2 : c2186 ? stack0_second2 : c2187 ? stack0_second31 : (c2361 || c2360) ? stack0_second36 : (c2188 && !c967) ? stack0_second2 : (c2157 && c1136) ? stack0_second2 : c2158 ? stack0_second2 : 'bz; */
            /* stack0_top50 <= (c2157 && c916) ? stack0_top2 : c2159 ? t947 : c2160 ? stack0_top2 : c2161 ? stack0_second2 : c2162 ? stack0_second2 : c2163 ? stack0_second2 : c2164 ? address0_top2 : c2246 ? stack0_top9 : c2247 ? stack0_second2 : c2166 ? stack0_top2 : c2167 ? stack0_top2 : c2168 ? stack0_second10 : c2169 ? stack0_second12 : c2170 ? stack0_second14 : c2171 ? stack0_second16 : c2172 ? stack0_top19 : c2173 ? stack0_second18 : c2174 ? stack0_top23 : c2175 ? stack0_top25 : c2176 ? stack0_top27 : (c2286 || c2284) ? stack0_top28 : c2178 ? stack0_top30 : c2179 ? stack0_top32 : c2180 ? stack0_top34 : c2181 ? stack0_top36 : c2182 ? stack0_top38 : c2212 ? stack0_second2 : (c2183 && !c964) ? stack0_top2 : c2184 ? stack0_top40 : c2185 ? stack0_top41 : c2186 ? stack0_top42 : c2187 ? stack0_second30 : (c2361 || c2360) ? stack0_top49 : (c2188 && !c967) ? stack0_top2 : (c2157 && c1136) ? stack0_top2 : c2158 ? stack0_top2 : 'bz; */
            t11 <= (c2157 && c916) ? t11 : c2159 ? t11 : c2160 ? t11 : c2161 ? t11 : c2162 ? t11 : c2163 ? t11 : c2164 ? t11 : c2246 ? t11 : c2247 ? t11 : c2166 ? t11 : c2167 ? t11 : c2168 ? t11 : c2169 ? t11 : c2170 ? t11 : c2171 ? t11 : c2172 ? t11 : c2173 ? t11 : c2174 ? stack0_top2 : c2175 ? stack0_top2 : c2176 ? stack0_top2 : (c2286 || c2284) ? t11 : c2178 ? stack0_top2 : c2179 ? stack0_top2 : c2180 ? stack0_top2 : c2181 ? stack0_top2 : c2182 ? stack0_top2 : c2212 ? t11 : (c2183 && !c964) ? t11 : c2184 ? t11 : c2185 ? t11 : c2186 ? stack0_top2 : c2187 ? t11 : (c2361 || c2360) ? t11 : (c2188 && !c967) ? t11 : (c2157 && c1136) ? t11 : c2158 ? t11 : 'bz;
            /* ip22 <= (ip21 + 1); */
            address0_pos2 <= address0_pos8;
            address0_second2 <= address0_second8;
            stack0_pos2 <= stack0_pos35;
            stack0_second2 <= stack0_second37;
            address0_top2 <= address0_top8;
            ip2 <= ip22;
            stack0_top2 <= stack0_top50;
            retro_main_state <= retro_main_L1_b198_S1;
          end
        end else begin
          _address_addr <= t843_inl7;
          _address_we <= 1;
          _address_req <= 1;
          _address_d <= address0_second2;
          memory_addr <= ip2;
          memory_we <= 0;
          memory_req <= 1;
          /* t843_inl7 <= (address0_pos2 - 2); */
          /* address0_pos7 <= (address0_pos2 + 1); */
          /* c2857 <= (c914 && !c915); */
          /* c2158 <= (c914 && !c915); */
          retro_main_state <= retro_main_L1_ifelse197_S1;
        end
      end
      retro_main_L1_ifelse197_S1: begin
        _address_req <= 0;
        /*wait for output of memory*/
        retro_main_state <= retro_main_L1_ifelse197_S2;
      end
      retro_main_L1_ifelse197_S2: begin
        t968 <= memory_q;
        memory_req <= 0;
        retro_main_state <= retro_main_L1_ifelse197_S3;
      end
      retro_main_L1_ifelse197_S3: begin
        /* ip20 <= (t968 - 1); */
        retro_main_state <= retro_main_L1_b198_S0;
      end
      retro_main_L1_ifthen11_S1: begin
        _stack_req <= 0;
        /*wait for output of memory*/
        retro_main_state <= retro_main_L1_ifthen11_S2;
      end
      retro_main_L1_ifthen11_S2: begin
        t947 <= memory_q;
        memory_req <= 0;
        retro_main_state <= retro_main_L1_b198_S0;
      end
      retro_main_L1_ifthen15_S1: begin
        _stack_req <= 0;
        retro_main_state <= retro_main_L1_b198_S0;
      end
      retro_main_L1_ifthen19_S1: begin
        /*wait for output of _stack*/
        retro_main_state <= retro_main_L1_ifthen19_S2;
      end
      retro_main_L1_ifthen19_S2: begin
        stack0_second5 <= _stack_q;
        _stack_req <= 0;
        retro_main_state <= retro_main_L1_b198_S0;
      end
      retro_main_L1_ifthen27_S1: begin
        /*wait for output of _stack*/
        _address_req <= 0;
        retro_main_state <= retro_main_L1_ifthen27_S2;
      end
      retro_main_L1_ifthen27_S2: begin
        stack0_second7 <= _stack_q;
        _stack_req <= 0;
        retro_main_state <= retro_main_L1_b198_S0;
      end
      retro_main_L1_ifthen31_S1: begin
        /*wait for output of _address*/
        _stack_req <= 0;
        retro_main_state <= retro_main_L1_ifthen31_S2;
      end
      retro_main_L1_ifthen31_S2: begin
        address0_second4 <= _address_q;
        _address_req <= 0;
        retro_main_state <= retro_main_L1_b198_S0;
      end
      retro_main_L1_ifthen44_S1: begin
        /*wait for output of memory*/
        retro_main_state <= retro_main_L1_ifthen44_S2;
      end
      retro_main_L1_ifthen44_S2: begin
        t954 <= memory_q;
        memory_req <= 0;
        retro_main_state <= retro_main_L1_ifthen44_S3;
      end
      retro_main_L1_ifthen44_S3: begin
        /* ip8 <= (t954 - 1); */
        retro_main_state <= retro_main_L1_b198_S0;
      end
      retro_main_L1_ifthen48_S1: begin
        /*wait for output of _address*/
        retro_main_state <= retro_main_L1_ifthen48_S2;
      end
      retro_main_L1_ifthen48_S2: begin
        address0_second5 <= _address_q;
        _address_req <= 0;
        retro_main_state <= retro_main_L1_b198_S0;
      end
      retro_main_L1_ifthen52_S1: begin
        _stack_addr <= t846_inl14;
        _stack_we <= 0;
        _stack_req <= 1;
        /*wait for output of _stack*/
        retro_main_state <= retro_main_L1_ifthen52_S2;
      end
      retro_main_L1_ifthen52_S2: begin
        /*wait for output of _stack*/
        stack0_second10 <= _stack_q;
        retro_main_state <= retro_main_L1_ifthen52_S3;
      end
      retro_main_L1_ifthen52_S3: begin
        stack0_second11 <= _stack_q;
        _stack_req <= 0;
        retro_main_state <= retro_main_L1_ifthen52_S4;
      end
      retro_main_L1_ifthen52_S4: begin
        if (c955) begin
          memory_addr <= ip10;
          memory_we <= 0;
          memory_req <= 1;
          /* c2890 <= (c2867 && c955); */
          retro_main_state <= retro_main_L1_ifthen55_S1;
        end else begin
          /* c2896 <= (c2867 && !c955); */
          /* t2660 <= c2277 ? ip11 : (c2168 && !c955) ? ip10 : 'bz; */
          retro_main_state <= retro_main_L1_b198_S0;
        end
      end
      retro_main_L1_ifthen61_S1: begin
        _stack_addr <= t846_inl16;
        _stack_we <= 0;
        _stack_req <= 1;
        /*wait for output of _stack*/
        retro_main_state <= retro_main_L1_ifthen61_S2;
      end
      retro_main_L1_ifthen61_S2: begin
        /*wait for output of _stack*/
        stack0_second12 <= _stack_q;
        retro_main_state <= retro_main_L1_ifthen61_S3;
      end
      retro_main_L1_ifthen61_S3: begin
        stack0_second13 <= _stack_q;
        _stack_req <= 0;
        retro_main_state <= retro_main_L1_ifthen61_S4;
      end
      retro_main_L1_ifthen61_S4: begin
        if (c957) begin
          memory_addr <= ip12;
          memory_we <= 0;
          memory_req <= 1;
          /* c2891 <= (c2868 && c957); */
          retro_main_state <= retro_main_L1_ifthen64_S1;
        end else begin
          /* c2897 <= (c2868 && !c957); */
          /* t2670 <= c2278 ? ip13 : (c2169 && !c957) ? ip12 : 'bz; */
          retro_main_state <= retro_main_L1_b198_S0;
        end
      end
      retro_main_L1_ifthen70_S1: begin
        _stack_addr <= t846_inl18;
        _stack_we <= 0;
        _stack_req <= 1;
        /*wait for output of _stack*/
        retro_main_state <= retro_main_L1_ifthen70_S2;
      end
      retro_main_L1_ifthen70_S2: begin
        /*wait for output of _stack*/
        stack0_second14 <= _stack_q;
        retro_main_state <= retro_main_L1_ifthen70_S3;
      end
      retro_main_L1_ifthen70_S3: begin
        stack0_second15 <= _stack_q;
        _stack_req <= 0;
        retro_main_state <= retro_main_L1_ifthen70_S4;
      end
      retro_main_L1_ifthen70_S4: begin
        if (c959) begin
          memory_addr <= ip14;
          memory_we <= 0;
          memory_req <= 1;
          /* c2892 <= (c2869 && c959); */
          retro_main_state <= retro_main_L1_ifthen73_S1;
        end else begin
          /* c2898 <= (c2869 && !c959); */
          /* t2680 <= c2279 ? ip15 : (c2170 && !c959) ? ip14 : 'bz; */
          retro_main_state <= retro_main_L1_b198_S0;
        end
      end
      retro_main_L1_ifthen79_S1: begin
        _stack_addr <= t846_inl20;
        _stack_we <= 0;
        _stack_req <= 1;
        /*wait for output of _stack*/
        retro_main_state <= retro_main_L1_ifthen79_S2;
      end
      retro_main_L1_ifthen79_S2: begin
        /*wait for output of _stack*/
        stack0_second16 <= _stack_q;
        retro_main_state <= retro_main_L1_ifthen79_S3;
      end
      retro_main_L1_ifthen79_S3: begin
        stack0_second17 <= _stack_q;
        _stack_req <= 0;
        retro_main_state <= retro_main_L1_ifthen79_S4;
      end
      retro_main_L1_ifthen79_S4: begin
        if (c961) begin
          memory_addr <= ip16;
          memory_we <= 0;
          memory_req <= 1;
          /* c2893 <= (c2870 && c961); */
          retro_main_state <= retro_main_L1_ifthen82_S1;
        end else begin
          /* c2899 <= (c2870 && !c961); */
          /* t2690 <= c2280 ? ip17 : (c2171 && !c961) ? ip16 : 'bz; */
          retro_main_state <= retro_main_L1_b198_S0;
        end
      end
      retro_main_L1_ifthen88_S1: begin
        /*wait for output of memory*/
        retro_main_state <= retro_main_L1_ifthen88_S2;
      end
      retro_main_L1_ifthen88_S2: begin
        stack0_top19 <= memory_q;
        memory_req <= 0;
        retro_main_state <= retro_main_L1_b198_S0;
      end
      retro_main_L1_ifthen92_S1: begin
        _stack_addr <= t846_inl22;
        _stack_we <= 0;
        _stack_req <= 1;
        /*wait for output of _stack*/
        memory_req <= 0;
        retro_main_state <= retro_main_L1_ifthen92_S2;
      end
      retro_main_L1_ifthen92_S2: begin
        /*wait for output of _stack*/
        stack0_second18 <= _stack_q;
        retro_main_state <= retro_main_L1_ifthen92_S3;
      end
      retro_main_L1_ifthen92_S3: begin
        stack0_second19 <= _stack_q;
        _stack_req <= 0;
        retro_main_state <= retro_main_L1_b198_S0;
      end
      retro_main_L1_ifthen96_S1: begin
        /*wait for output of _stack*/
        retro_main_state <= retro_main_L1_ifthen96_S2;
      end
      retro_main_L1_ifthen96_S2: begin
        stack0_second20 <= _stack_q;
        _stack_req <= 0;
        retro_main_state <= retro_main_L1_b198_S0;
      end
      retro_main_L1_ifthen100_S1: begin
        /*wait for output of _stack*/
        retro_main_state <= retro_main_L1_ifthen100_S2;
      end
      retro_main_L1_ifthen100_S2: begin
        stack0_second21 <= _stack_q;
        _stack_req <= 0;
        retro_main_state <= retro_main_L1_b198_S0;
      end
      retro_main_L1_ifthen104_S1: begin
        /*wait for output of _stack*/
        retro_main_state <= retro_main_L1_ifthen104_S2;
      end
      retro_main_L1_ifthen104_S2: begin
        stack0_second22 <= _stack_q;
        _stack_req <= 0;
        retro_main_state <= retro_main_L1_b198_S0;
      end
      retro_main_L1_ifthen112_S1: begin
        /*wait for output of _stack*/
        retro_main_state <= retro_main_L1_ifthen112_S2;
      end
      retro_main_L1_ifthen112_S2: begin
        stack0_second24 <= _stack_q;
        _stack_req <= 0;
        retro_main_state <= retro_main_L1_b198_S0;
      end
      retro_main_L1_ifthen116_S1: begin
        /*wait for output of _stack*/
        retro_main_state <= retro_main_L1_ifthen116_S2;
      end
      retro_main_L1_ifthen116_S2: begin
        stack0_second25 <= _stack_q;
        _stack_req <= 0;
        retro_main_state <= retro_main_L1_b198_S0;
      end
      retro_main_L1_ifthen120_S1: begin
        /*wait for output of _stack*/
        retro_main_state <= retro_main_L1_ifthen120_S2;
      end
      retro_main_L1_ifthen120_S2: begin
        stack0_second26 <= _stack_q;
        _stack_req <= 0;
        retro_main_state <= retro_main_L1_b198_S0;
      end
      retro_main_L1_ifthen124_S1: begin
        /*wait for output of _stack*/
        retro_main_state <= retro_main_L1_ifthen124_S2;
      end
      retro_main_L1_ifthen124_S2: begin
        stack0_second27 <= _stack_q;
        _stack_req <= 0;
        retro_main_state <= retro_main_L1_b198_S0;
      end
      retro_main_L1_ifthen128_S1: begin
        /*wait for output of _stack*/
        retro_main_state <= retro_main_L1_ifthen128_S2;
      end
      retro_main_L1_ifthen128_S2: begin
        stack0_second28 <= _stack_q;
        _stack_req <= 0;
        retro_main_state <= retro_main_L1_b198_S0;
      end
      retro_main_L1_ifthen153_S1: begin
        _stack_addr <= t846_inl34;
        _stack_we <= 0;
        _stack_req <= 1;
        /*wait for output of _stack*/
        retro_main_state <= retro_main_L1_ifthen153_S2;
      end
      retro_main_L1_ifthen153_S2: begin
        /*wait for output of _stack*/
        stack0_second30 <= _stack_q;
        retro_main_state <= retro_main_L1_ifthen153_S3;
      end
      retro_main_L1_ifthen153_S3: begin
        stack0_second31 <= _stack_q;
        _stack_req <= 0;
        retro_main_state <= retro_main_L1_b198_S0;
      end
      retro_main_L1_ifthen157_S1: begin
        /* c967 <= (t966 == 0); */
        if (c967) begin
          array998[0] <= 1;
          t847_inl51 <= array998[1];
          /* c2895 <= (c2887 && c967); */
          /* c2217 <= (c2188 && c967); */
          retro_main_state <= retro_main_L1_ifthen160_S1;
        end else begin
          a6 <= (c2157 && c916) ? a6 : c2159 ? a6 : c2160 ? a6 : c2161 ? a6 : c2162 ? a6 : c2163 ? a6 : c2164 ? a6 : c2246 ? a6 : c2247 ? a6 : c2166 ? a6 : c2167 ? a6 : c2168 ? stack0_top2 : c2169 ? stack0_top2 : c2170 ? stack0_top2 : c2171 ? stack0_top2 : c2172 ? a6 : c2173 ? a6 : c2174 ? a6 : c2175 ? a6 : c2176 ? a6 : (c2286 || c2284) ? a6 : c2178 ? a6 : c2179 ? a6 : c2180 ? a6 : c2181 ? a6 : c2182 ? a6 : c2212 ? a6 : (c2183 && !c964) ? a6 : c2184 ? a6 : c2185 ? a6 : c2186 ? a6 : c2187 ? a6 : (c2361 || c2360) ? a6 : (c2188 && !c967) ? a6 : (c2157 && c1136) ? a6 : c2158 ? a6 : 'bz;
          /* address0_pos8 <= (c2157 && c916) ? address0_pos2 : c2159 ? address0_pos2 : c2160 ? address0_pos2 : c2161 ? address0_pos2 : c2162 ? address0_pos2 : c2163 ? address0_pos3 : c2164 ? address0_pos4 : c2246 ? address0_pos2 : c2247 ? address0_pos2 : c2166 ? address0_pos2 : c2167 ? address0_pos5 : c2168 ? address0_pos2 : c2169 ? address0_pos2 : c2170 ? address0_pos2 : c2171 ? address0_pos2 : c2172 ? address0_pos2 : c2173 ? address0_pos2 : c2174 ? address0_pos2 : c2175 ? address0_pos2 : c2176 ? address0_pos2 : (c2286 || c2284) ? address0_pos2 : c2178 ? address0_pos2 : c2179 ? address0_pos2 : c2180 ? address0_pos2 : c2181 ? address0_pos2 : c2182 ? address0_pos2 : c2212 ? address0_pos6 : (c2183 && !c964) ? address0_pos2 : c2184 ? address0_pos2 : c2185 ? address0_pos2 : c2186 ? address0_pos2 : c2187 ? address0_pos2 : (c2361 || c2360) ? address0_pos2 : (c2188 && !c967) ? address0_pos2 : (c2157 && c1136) ? address0_pos2 : c2158 ? address0_pos7 : 'bz; */
          /* address0_second8 <= (c2157 && c916) ? address0_second2 : c2159 ? address0_second2 : c2160 ? address0_second2 : c2161 ? address0_second2 : c2162 ? address0_second2 : c2163 ? address0_top2 : c2164 ? address0_second4 : c2246 ? address0_second2 : c2247 ? address0_second2 : c2166 ? address0_second2 : c2167 ? address0_second5 : c2168 ? address0_second2 : c2169 ? address0_second2 : c2170 ? address0_second2 : c2171 ? address0_second2 : c2172 ? address0_second2 : c2173 ? address0_second2 : c2174 ? address0_second2 : c2175 ? address0_second2 : c2176 ? address0_second2 : (c2286 || c2284) ? address0_second2 : c2178 ? address0_second2 : c2179 ? address0_second2 : c2180 ? address0_second2 : c2181 ? address0_second2 : c2182 ? address0_second2 : c2212 ? address0_second6 : (c2183 && !c964) ? address0_second2 : c2184 ? address0_second2 : c2185 ? address0_second2 : c2186 ? address0_second2 : c2187 ? address0_second2 : (c2361 || c2360) ? address0_second2 : (c2188 && !c967) ? address0_second2 : (c2157 && c1136) ? address0_second2 : c2158 ? address0_top2 : 'bz; */
          /* address0_top8 <= (c2157 && c916) ? address0_top2 : c2159 ? address0_top2 : c2160 ? address0_top2 : c2161 ? address0_top2 : c2162 ? address0_top2 : c2163 ? stack0_top2 : c2164 ? address0_second2 : c2246 ? address0_top2 : c2247 ? address0_top2 : c2166 ? address0_top2 : c2167 ? address0_second2 : c2168 ? address0_top2 : c2169 ? address0_top2 : c2170 ? address0_top2 : c2171 ? address0_top2 : c2172 ? address0_top2 : c2173 ? address0_top2 : c2174 ? address0_top2 : c2175 ? address0_top2 : c2176 ? address0_top2 : (c2286 || c2284) ? address0_top2 : c2178 ? address0_top2 : c2179 ? address0_top2 : c2180 ? address0_top2 : c2181 ? address0_top2 : c2182 ? address0_top2 : c2212 ? address0_second2 : (c2183 && !c964) ? address0_top2 : c2184 ? address0_top2 : c2185 ? address0_top2 : c2186 ? address0_top2 : c2187 ? address0_top2 : (c2361 || c2360) ? address0_top2 : (c2188 && !c967) ? address0_top2 : (c2157 && c1136) ? address0_top2 : c2158 ? ip2 : 'bz; */
          b6 <= (c2157 && c916) ? b6 : c2159 ? b6 : c2160 ? b6 : c2161 ? b6 : c2162 ? b6 : c2163 ? b6 : c2164 ? b6 : c2246 ? b6 : c2247 ? b6 : c2166 ? b6 : c2167 ? b6 : c2168 ? stack0_second2 : c2169 ? stack0_second2 : c2170 ? stack0_second2 : c2171 ? stack0_second2 : c2172 ? b6 : c2173 ? b6 : c2174 ? b6 : c2175 ? b6 : c2176 ? b6 : (c2286 || c2284) ? b6 : c2178 ? b6 : c2179 ? b6 : c2180 ? b6 : c2181 ? b6 : c2182 ? b6 : c2212 ? b6 : (c2183 && !c964) ? b6 : c2184 ? b6 : c2185 ? b6 : c2186 ? b6 : c2187 ? b6 : (c2361 || c2360) ? b6 : (c2188 && !c967) ? b6 : (c2157 && c1136) ? b6 : c2158 ? b6 : 'bz;
          /* ip21 <= (c2157 && c916) ? ip2 : c2159 ? ip3 : c2160 ? ip2 : c2161 ? ip2 : c2162 ? ip2 : c2163 ? ip2 : c2164 ? ip2 : c2246 ? ip5 : c2247 ? ip6 : c2166 ? ip8 : c2167 ? address0_top2 : c2168 ? t2660 : c2169 ? t2670 : c2170 ? t2680 : c2171 ? t2690 : c2172 ? ip2 : c2173 ? ip2 : c2174 ? ip2 : c2175 ? ip2 : c2176 ? ip2 : (c2286 || c2284) ? ip2 : c2178 ? ip2 : c2179 ? ip2 : c2180 ? ip2 : c2181 ? ip2 : c2182 ? ip2 : c2212 ? address0_top2 : (c2183 && !c964) ? ip2 : c2184 ? ip2 : c2185 ? ip2 : c2186 ? ip2 : c2187 ? ip2 : (c2361 || c2360) ? ip_inl514 : (c2188 && !c967) ? ip2 : (c2157 && c1136) ? ip2 : c2158 ? ip20 : 'bz; */
          /* stack0_pos35 <= (c2157 && c916) ? stack0_pos2 : c2159 ? stack0_pos3 : c2160 ? stack0_pos4 : c2161 ? stack0_pos5 : c2162 ? stack0_pos2 : c2163 ? stack0_pos6 : c2164 ? stack0_pos7 : c2246 ? stack0_pos2 : c2247 ? stack0_pos8 : c2166 ? stack0_pos2 : c2167 ? stack0_pos2 : c2168 ? stack0_pos10 : c2169 ? stack0_pos12 : c2170 ? stack0_pos14 : c2171 ? stack0_pos16 : c2172 ? stack0_pos2 : c2173 ? stack0_pos18 : c2174 ? stack0_pos19 : c2175 ? stack0_pos20 : c2176 ? stack0_pos21 : (c2286 || c2284) ? stack0_pos2 : c2178 ? stack0_pos22 : c2179 ? stack0_pos23 : c2180 ? stack0_pos24 : c2181 ? stack0_pos25 : c2182 ? stack0_pos26 : c2212 ? stack0_pos27 : (c2183 && !c964) ? stack0_pos2 : c2184 ? stack0_pos2 : c2185 ? stack0_pos2 : c2186 ? stack0_pos2 : c2187 ? stack0_pos29 : (c2361 || c2360) ? stack0_pos34 : (c2188 && !c967) ? stack0_pos2 : (c2157 && c1136) ? stack0_pos2 : c2158 ? stack0_pos2 : 'bz; */
          /* stack0_second37 <= (c2157 && c916) ? stack0_second2 : c2159 ? stack0_top2 : c2160 ? stack0_top2 : c2161 ? stack0_second5 : c2162 ? stack0_top2 : c2163 ? stack0_second7 : c2164 ? stack0_top2 : c2246 ? stack0_second2 : c2247 ? stack0_second9 : c2166 ? stack0_second2 : c2167 ? stack0_second2 : c2168 ? stack0_second11 : c2169 ? stack0_second13 : c2170 ? stack0_second15 : c2171 ? stack0_second17 : c2172 ? stack0_second2 : c2173 ? stack0_second19 : c2174 ? stack0_second20 : c2175 ? stack0_second21 : c2176 ? stack0_second22 : (c2286 || c2284) ? stack0_second23 : c2178 ? stack0_second24 : c2179 ? stack0_second25 : c2180 ? stack0_second26 : c2181 ? stack0_second27 : c2182 ? stack0_second28 : c2212 ? stack0_second29 : (c2183 && !c964) ? stack0_second2 : c2184 ? stack0_second2 : c2185 ? stack0_second2 : c2186 ? stack0_second2 : c2187 ? stack0_second31 : (c2361 || c2360) ? stack0_second36 : (c2188 && !c967) ? stack0_second2 : (c2157 && c1136) ? stack0_second2 : c2158 ? stack0_second2 : 'bz; */
          /* stack0_top50 <= (c2157 && c916) ? stack0_top2 : c2159 ? t947 : c2160 ? stack0_top2 : c2161 ? stack0_second2 : c2162 ? stack0_second2 : c2163 ? stack0_second2 : c2164 ? address0_top2 : c2246 ? stack0_top9 : c2247 ? stack0_second2 : c2166 ? stack0_top2 : c2167 ? stack0_top2 : c2168 ? stack0_second10 : c2169 ? stack0_second12 : c2170 ? stack0_second14 : c2171 ? stack0_second16 : c2172 ? stack0_top19 : c2173 ? stack0_second18 : c2174 ? stack0_top23 : c2175 ? stack0_top25 : c2176 ? stack0_top27 : (c2286 || c2284) ? stack0_top28 : c2178 ? stack0_top30 : c2179 ? stack0_top32 : c2180 ? stack0_top34 : c2181 ? stack0_top36 : c2182 ? stack0_top38 : c2212 ? stack0_second2 : (c2183 && !c964) ? stack0_top2 : c2184 ? stack0_top40 : c2185 ? stack0_top41 : c2186 ? stack0_top42 : c2187 ? stack0_second30 : (c2361 || c2360) ? stack0_top49 : (c2188 && !c967) ? stack0_top2 : (c2157 && c1136) ? stack0_top2 : c2158 ? stack0_top2 : 'bz; */
          t11 <= (c2157 && c916) ? t11 : c2159 ? t11 : c2160 ? t11 : c2161 ? t11 : c2162 ? t11 : c2163 ? t11 : c2164 ? t11 : c2246 ? t11 : c2247 ? t11 : c2166 ? t11 : c2167 ? t11 : c2168 ? t11 : c2169 ? t11 : c2170 ? t11 : c2171 ? t11 : c2172 ? t11 : c2173 ? t11 : c2174 ? stack0_top2 : c2175 ? stack0_top2 : c2176 ? stack0_top2 : (c2286 || c2284) ? t11 : c2178 ? stack0_top2 : c2179 ? stack0_top2 : c2180 ? stack0_top2 : c2181 ? stack0_top2 : c2182 ? stack0_top2 : c2212 ? t11 : (c2183 && !c964) ? t11 : c2184 ? t11 : c2185 ? t11 : c2186 ? stack0_top2 : c2187 ? t11 : (c2361 || c2360) ? t11 : (c2188 && !c967) ? t11 : (c2157 && c1136) ? t11 : c2158 ? t11 : 'bz;
          /* ip22 <= (ip21 + 1); */
          address0_pos2 <= address0_pos8;
          address0_second2 <= address0_second8;
          stack0_pos2 <= stack0_pos35;
          stack0_second2 <= stack0_second37;
          address0_top2 <= address0_top8;
          ip2 <= ip22;
          stack0_top2 <= stack0_top50;
          retro_main_state <= retro_main_L1_b198_S1;
        end
      end
      retro_main_L1_ifthen38_S1: begin
        /*wait for output of memory*/
        retro_main_state <= retro_main_L1_ifthen38_S2;
      end
      retro_main_L1_ifthen38_S2: begin
        t953 <= memory_q;
        memory_req <= 0;
        retro_main_state <= retro_main_L1_ifthen38_S3;
      end
      retro_main_L1_ifthen38_S3: begin
        /* ip5 <= (t953 - 1); */
        retro_main_state <= retro_main_L1_b198_S0;
      end
      retro_main_L1_ifelse41_S1: begin
        /*wait for output of _stack*/
        retro_main_state <= retro_main_L1_ifelse41_S2;
      end
      retro_main_L1_ifelse41_S2: begin
        stack0_second9 <= _stack_q;
        _stack_req <= 0;
        retro_main_state <= retro_main_L1_b198_S0;
      end
      retro_main_L1_ifthen55_S1: begin
        /*wait for output of memory*/
        retro_main_state <= retro_main_L1_ifthen55_S2;
      end
      retro_main_L1_ifthen55_S2: begin
        t956 <= memory_q;
        memory_req <= 0;
        retro_main_state <= retro_main_L1_ifthen55_S3;
      end
      retro_main_L1_ifthen55_S3: begin
        /* ip11 <= (t956 - 1); */
        retro_main_state <= retro_main_L1_b603_S0;
      end
      retro_main_L1_ifthen64_S1: begin
        /*wait for output of memory*/
        retro_main_state <= retro_main_L1_ifthen64_S2;
      end
      retro_main_L1_ifthen64_S2: begin
        t958 <= memory_q;
        memory_req <= 0;
        retro_main_state <= retro_main_L1_ifthen64_S3;
      end
      retro_main_L1_ifthen64_S3: begin
        /* ip13 <= (t958 - 1); */
        retro_main_state <= retro_main_L1_b604_S0;
      end
      retro_main_L1_ifthen73_S1: begin
        /*wait for output of memory*/
        retro_main_state <= retro_main_L1_ifthen73_S2;
      end
      retro_main_L1_ifthen73_S2: begin
        t960 <= memory_q;
        memory_req <= 0;
        retro_main_state <= retro_main_L1_ifthen73_S3;
      end
      retro_main_L1_ifthen73_S3: begin
        /* ip15 <= (t960 - 1); */
        retro_main_state <= retro_main_L1_b605_S0;
      end
      retro_main_L1_ifthen82_S1: begin
        /*wait for output of memory*/
        retro_main_state <= retro_main_L1_ifthen82_S2;
      end
      retro_main_L1_ifthen82_S2: begin
        t962 <= memory_q;
        memory_req <= 0;
        retro_main_state <= retro_main_L1_ifthen82_S3;
      end
      retro_main_L1_ifthen82_S3: begin
        /* ip17 <= (t962 - 1); */
        retro_main_state <= retro_main_L1_b606_S0;
      end
      retro_main_L1_ifthen135_S1: begin
        /*wait for output of _address*/
        /*wait for output of _stack*/
        retro_main_state <= retro_main_L1_ifthen135_S2;
      end
      retro_main_L1_ifthen135_S2: begin
        address0_second6 <= _address_q;
        _address_req <= 0;
        stack0_second29 <= _stack_q;
        _stack_req <= 0;
        retro_main_state <= retro_main_L1_b198_S0;
      end
      retro_main_L1_ifthen160_S1: begin
        /* c848_inl51 <= (t847_inl51 == 1); */
        if (c848_inl51) begin
          /* c2901 <= (c2895 && c848_inl51); */
          /* c2243 <= (c2217 && c848_inl51); */
          retro_main_state <= retro_main_L2_while427_S0;
        end else begin
          t852_inl51 <= array998[2];
          /* c2914 <= (c2895 && !c848_inl51); */
          /* c2290 <= (c2217 && !c848_inl51); */
          /* c2915 <= (c2901 && !c851_inl51); */
          /* c2291 <= (c2243 && !c851_inl51); */
          retro_main_state <= retro_main_L1_b443_S1;
        end
      end
      retro_main_L1_b603_S0: begin
        /* c2896 <= (c2867 && !c955); */
        /* t2660 <= c2277 ? ip11 : (c2168 && !c955) ? ip10 : 'bz; */
        retro_main_state <= retro_main_L1_b198_S0;
      end
      retro_main_L1_b604_S0: begin
        /* c2897 <= (c2868 && !c957); */
        /* t2670 <= c2278 ? ip13 : (c2169 && !c957) ? ip12 : 'bz; */
        retro_main_state <= retro_main_L1_b198_S0;
      end
      retro_main_L1_b605_S0: begin
        /* c2898 <= (c2869 && !c959); */
        /* t2680 <= c2279 ? ip15 : (c2170 && !c959) ? ip14 : 'bz; */
        retro_main_state <= retro_main_L1_b198_S0;
      end
      retro_main_L1_b606_S0: begin
        /* c2899 <= (c2870 && !c961); */
        /* t2690 <= c2280 ? ip17 : (c2171 && !c961) ? ip16 : 'bz; */
        retro_main_state <= retro_main_L1_b198_S0;
      end
      retro_main_L1_exit396_S0: begin
        i_inl2_inl493 <= 0;
        n_inl2_inl493 <= 0;
        test_bit_inl2_inl493 <= 1073741824;
        /* x_inl2_inl49 <= abs_b_inl492; */
        /* c2904 <= (c2876 && !c986_inl1_inl49); */
        retro_main_state <= retro_main_L1_exit396_S1;
      end
      retro_main_L1_exit396_S1: begin
        retro_main_state <= retro_main_L21_fortest399_S0;
      end
      retro_main_L1_whileexit429_S1: begin
        io_ports_req <= 0;
        retro_main_state <= retro_main_L3_while432_S0;
      end
      retro_main_L1_whileexit434_S1: begin
        io_ports_addr <= 1;
        io_ports_we <= 1;
        io_ports_req <= 1;
        io_ports_d <= 0;
        /*wait for output of io_ports*/
        retro_main_state <= retro_main_L1_whileexit434_S2;
      end
      retro_main_L1_whileexit434_S2: begin
        io_ports_req <= 0;
        char_c_inl1_inl51 <= io_ports_q;
        retro_main_state <= retro_main_L4_while437_S0;
      end
      retro_main_L1_exit402_S0: begin
        c_bit_inl493 <= 0;
        i_inl493 <= 0;
        abs_a_inl493 <= abs_a_inl492;
        /* find_zero_len_result2_inl494 <= c2284 ? n_inl2_inl493 : (c2177 || c2256) ? 0 : 'bz; */
        /* c2286 <= (c2177 || c2256); */
        /* c2910 <= ((c2904 || c2902) && !c986_inl2_inl49); */
        /* abs_b_inl493 <= (abs_b_inl492 << find_zero_len_result2_inl494); */
        /* t486_inl49 <= (find_zero_len_result2_inl494 + 1); */
        abs_b_inl494 <= abs_b_inl493;
        retro_main_state <= retro_main_L1_exit402_S1;
      end
      retro_main_L1_exit402_S1: begin
        retro_main_state <= retro_main_L22_fortest404_S0;
      end
      retro_main_L1_whileexit439_S1: begin
        t850_inl51 <= array998[1];
        retro_main_state <= retro_main_L1_whileexit439_S2;
      end
      retro_main_L1_whileexit439_S2: begin
        /* c851_inl51 <= (t850_inl51 == 13); */
        /* c2288 <= (c2243 && c851_inl51); */
        if (c851_inl51) begin
          array998[1] <= 10;
          /* c2912 <= (c2901 && c851_inl51); */
          retro_main_state <= retro_main_L1_b443_S0;
        end else begin
          t852_inl51 <= array998[2];
          /* c2914 <= (c2895 && !c848_inl51); */
          /* c2290 <= (c2217 && !c848_inl51); */
          /* c2915 <= (c2901 && !c851_inl51); */
          /* c2291 <= (c2243 && !c851_inl51); */
          retro_main_state <= retro_main_L1_b443_S1;
        end
      end
      retro_main_L1_forelse409_S2: begin
        /* stack0_top28 <= retro_divmod_result492[0]; */
        /* stack0_second23 <= retro_divmod_result492[1]; */
        retro_main_state <= retro_main_L1_b198_S0;
      end
      retro_main_L1_b443_S0: begin
        t852_inl51 <= array998[2];
        /* c2914 <= (c2895 && !c848_inl51); */
        /* c2290 <= (c2217 && !c848_inl51); */
        /* c2915 <= (c2901 && !c851_inl51); */
        /* c2291 <= (c2243 && !c851_inl51); */
        retro_main_state <= retro_main_L1_b443_S1;
      end
      retro_main_L1_b443_S1: begin
        /* c853_inl51 <= (t852_inl51 == 1); */
        if (c853_inl51) begin
          /* c854_inl51 <= (stack0_top2 > 0); */
          /* c855_inl51 <= (stack0_top2 < 128); */
          /* c856_inl51 <= (c854_inl51 && c855_inl51); */
          /* c2916 <= (((c2914 || c2915) || c2912) && c853_inl51); */
          /* c2295 <= (((c2290 || c2291) || c2288) && c853_inl51); */
          if (c856_inl51) begin
            /* c857_inl51 <= (stack0_top2 == 8); */
            /* c2917 <= (c2916 && c856_inl51); */
            /* c2297 <= (c2295 && c856_inl51); */
            if (c857_inl51) begin
              _stack_addr <= t846_inl2_inl51;
              _stack_we <= 0;
              _stack_req <= 1;
              /* stack0_pos30 <= (stack0_pos2 - 1); */
              /* t846_inl2_inl51 <= (stack0_pos30 - 2); */
              /* c2919 <= (c2917 && c857_inl51); */
              /* c2300 <= (c2297 && c857_inl51); */
              retro_main_state <= retro_main_L1_ifthen446_S1;
            end else begin
              _stack_addr <= t846_inl3_inl51;
              _stack_we <= 0;
              _stack_req <= 1;
              /* stack0_pos31 <= (stack0_pos2 - 1); */
              /* t846_inl3_inl51 <= (stack0_pos31 - 2); */
              /* c2920 <= (c2917 && !c857_inl51); */
              /* c2301 <= (c2297 && !c857_inl51); */
              retro_main_state <= retro_main_L1_ifelse569_S1;
            end
          end else begin
            _stack_addr <= t846_inl4_inl51;
            _stack_we <= 0;
            _stack_req <= 1;
            /* stack0_pos32 <= (stack0_pos2 - 1); */
            /* t846_inl4_inl51 <= (stack0_pos32 - 2); */
            /* c2918 <= (c2916 && !c856_inl51); */
            /* c2298 <= (c2295 && !c856_inl51); */
            retro_main_state <= retro_main_L1_ifelse594_S1;
          end
        end else begin
          t859_inl51 <= array998[4];
          /* c2938 <= (((c2914 || c2915) || c2912) && !c853_inl51); */
          /* c2328 <= (((c2290 || c2291) || c2288) && !c853_inl51); */
          /* c2939 <= ((c2918 || c2932) || c2933); */
          /* stack0_pos34 <= ((c2298 || c2322) || c2323) ? stack0_pos33 : (((c2290 || c2291) || c2288) && !c853_inl51) ? stack0_pos2 : 'bz; */
          /* stack0_second36 <= ((c2298 || c2322) || c2323) ? stack0_second35 : (((c2290 || c2291) || c2288) && !c853_inl51) ? stack0_second2 : 'bz; */
          /* stack0_top49 <= ((c2298 || c2322) || c2323) ? stack0_second2 : (((c2290 || c2291) || c2288) && !c853_inl51) ? stack0_top2 : 'bz; */
          /* c2329 <= ((c2298 || c2322) || c2323); */
          retro_main_state <= retro_main_L1_b520_S1;
        end
      end
      retro_main_L1_ifelse594_S1: begin
        /*wait for output of _stack*/
        retro_main_state <= retro_main_L1_ifelse594_S2;
      end
      retro_main_L1_ifelse594_S2: begin
        stack0_second34 <= _stack_q;
        _stack_req <= 0;
        retro_main_state <= retro_main_L1_b502_S0;
      end
      retro_main_L1_ifthen446_S1: begin
        /*wait for output of _stack*/
        retro_main_state <= retro_main_L1_ifthen446_S2;
      end
      retro_main_L1_ifthen446_S2: begin
        stack0_second32 <= _stack_q;
        _stack_req <= 0;
        retro_main_state <= retro_main_L8_while453_S0;
      end
      retro_main_L1_ifelse569_S1: begin
        /*wait for output of _stack*/
        retro_main_state <= retro_main_L1_ifelse569_S2;
      end
      retro_main_L1_ifelse569_S2: begin
        stack0_second33 <= _stack_q;
        _stack_req <= 0;
        retro_main_state <= retro_main_L5_while576_S0;
      end
      retro_main_L1_whileexit455_S1: begin
        io_ports_addr <= 1;
        io_ports_we <= 1;
        io_ports_req <= 1;
        io_ports_d <= 1;
        retro_main_state <= retro_main_L1_whileexit455_S2;
      end
      retro_main_L1_whileexit455_S2: begin
        io_ports_req <= 0;
        retro_main_state <= retro_main_L9_while458_S0;
      end
      retro_main_L1_whileexit578_S1: begin
        io_ports_addr <= 1;
        io_ports_we <= 1;
        io_ports_req <= 1;
        io_ports_d <= 1;
        retro_main_state <= retro_main_L1_whileexit578_S2;
      end
      retro_main_L1_whileexit578_S2: begin
        io_ports_req <= 0;
        retro_main_state <= retro_main_L6_while581_S0;
      end
      retro_main_L1_whileexit460_S1: begin
        io_ports_req <= 0;
        retro_main_state <= retro_main_L10_while463_S0;
      end
      retro_main_L1_whileexit583_S1: begin
        io_ports_req <= 0;
        retro_main_state <= retro_main_L7_while586_S0;
      end
      retro_main_L1_whileexit472_S1: begin
        io_ports_addr <= 1;
        io_ports_we <= 1;
        io_ports_req <= 1;
        io_ports_d <= 1;
        retro_main_state <= retro_main_L1_whileexit472_S2;
      end
      retro_main_L1_whileexit472_S2: begin
        io_ports_req <= 0;
        retro_main_state <= retro_main_L12_while475_S0;
      end
      retro_main_L1_whileexit477_S1: begin
        io_ports_req <= 0;
        retro_main_state <= retro_main_L13_while480_S0;
      end
      retro_main_L1_whileexit489_S1: begin
        io_ports_addr <= 1;
        io_ports_we <= 1;
        io_ports_req <= 1;
        io_ports_d <= 1;
        retro_main_state <= retro_main_L1_whileexit489_S2;
      end
      retro_main_L1_whileexit489_S2: begin
        io_ports_req <= 0;
        retro_main_state <= retro_main_L15_while492_S0;
      end
      retro_main_L1_whileexit494_S1: begin
        io_ports_req <= 0;
        retro_main_state <= retro_main_L16_while497_S0;
      end
      retro_main_L1_b502_S0: begin
        /* stack0_pos33 <= (c2300 && c985_inl3_inl7_inl51) ? stack0_pos30 : (c2301 && c985_inl3_inl8_inl51) ? stack0_pos31 : c2298 ? stack0_pos32 : 'bz; */
        /* c2932 <= (c2920 && c985_inl3_inl8_inl51); */
        /* c2933 <= (c2919 && c985_inl3_inl7_inl51); */
        /* stack0_second35 <= (c2300 && c985_inl3_inl7_inl51) ? stack0_second32 : (c2301 && c985_inl3_inl8_inl51) ? stack0_second33 : c2298 ? stack0_second34 : 'bz; */
        /* c2322 <= (c2301 && c985_inl3_inl8_inl51); */
        /* c2323 <= (c2300 && c985_inl3_inl7_inl51); */
        retro_main_state <= retro_main_L17_while505_S0;
      end
      retro_main_L1_whileexit507_S1: begin
        io_ports_req <= 0;
        retro_main_state <= retro_main_L18_while510_S0;
      end
      retro_main_L1_whileexit512_S1: begin
        io_ports_req <= 0;
        retro_main_state <= retro_main_L19_while515_S0;
      end
      retro_main_L1_b520_S0: begin
        t859_inl51 <= array998[4];
        /* c2938 <= (((c2914 || c2915) || c2912) && !c853_inl51); */
        /* c2328 <= (((c2290 || c2291) || c2288) && !c853_inl51); */
        /* c2939 <= ((c2918 || c2932) || c2933); */
        /* stack0_pos34 <= ((c2298 || c2322) || c2323) ? stack0_pos33 : (((c2290 || c2291) || c2288) && !c853_inl51) ? stack0_pos2 : 'bz; */
        /* stack0_second36 <= ((c2298 || c2322) || c2323) ? stack0_second35 : (((c2290 || c2291) || c2288) && !c853_inl51) ? stack0_second2 : 'bz; */
        /* stack0_top49 <= ((c2298 || c2322) || c2323) ? stack0_second2 : (((c2290 || c2291) || c2288) && !c853_inl51) ? stack0_top2 : 'bz; */
        /* c2329 <= ((c2298 || c2322) || c2323); */
        retro_main_state <= retro_main_L1_b520_S1;
      end
      retro_main_L1_b520_S1: begin
        /* c860_inl51 <= (t859_inl51 == 1); */
        /* c2330 <= ((c2328 || c2329) && c860_inl51); */
        if (c860_inl51) begin
          array998[4] <= 0;
          /* c2940 <= ((c2938 || c2939) && c860_inl51); */
          retro_main_state <= retro_main_L1_b522_S0;
        end else begin
          t861_inl51 <= array998[4];
          /* c2941 <= ((c2938 || c2939) && !c860_inl51); */
          /* c2331 <= ((c2328 || c2329) && !c860_inl51); */
          retro_main_state <= retro_main_L1_b522_S1;
        end
      end
      retro_main_L1_b522_S0: begin
        t861_inl51 <= array998[4];
        /* c2941 <= ((c2938 || c2939) && !c860_inl51); */
        /* c2331 <= ((c2328 || c2329) && !c860_inl51); */
        retro_main_state <= retro_main_L1_b522_S1;
      end
      retro_main_L1_b522_S1: begin
        /* c862_inl51 <= (t861_inl51 == 2); */
        /* c2332 <= ((c2331 || c2330) && c862_inl51); */
        if (c862_inl51) begin
          array998[4] <= 0;
          /* c2942 <= ((c2941 || c2940) && c862_inl51); */
          retro_main_state <= retro_main_L1_b524_S0;
        end else begin
          t863_inl51 <= array998[4];
          t865_inl51 <= array998[4];
          t867_inl51 <= array998[4];
          t869_inl51 <= array998[4];
          t871_inl51 <= array998[4];
          t873_inl51 <= array998[4];
          t875_inl51 <= array998[4];
          /* c2943 <= ((c2941 || c2940) && !c862_inl51); */
          /* c2333 <= ((c2331 || c2330) && !c862_inl51); */
          retro_main_state <= retro_main_L1_b524_S1;
        end
      end
      retro_main_L1_b524_S0: begin
        t863_inl51 <= array998[4];
        t865_inl51 <= array998[4];
        t867_inl51 <= array998[4];
        t869_inl51 <= array998[4];
        t871_inl51 <= array998[4];
        t873_inl51 <= array998[4];
        t875_inl51 <= array998[4];
        /* c2943 <= ((c2941 || c2940) && !c862_inl51); */
        /* c2333 <= ((c2331 || c2330) && !c862_inl51); */
        retro_main_state <= retro_main_L1_b524_S1;
      end
      retro_main_L1_b524_S1: begin
        /* c864_inl51 <= (t863_inl51 == -1); */
        /* c866_inl51 <= (t865_inl51 == -2); */
        /* c868_inl51 <= (t867_inl51 == -3); */
        /* c870_inl51 <= (t869_inl51 == -4); */
        /* c872_inl51 <= (t871_inl51 == -5); */
        /* c874_inl51 <= (t873_inl51 == -6); */
        /* c876_inl51 <= (t875_inl51 == -7); */
        /* c1084_inl51 <= (!c864_inl51 && c866_inl51); */
        /* c1085_inl51 <= ((!c864_inl51 && !c866_inl51) && c868_inl51); */
        /* c1086_inl51 <= (((!c864_inl51 && !c866_inl51) && !c868_inl51) && c870_inl51); */
        /* c1087_inl51 <= ((((!c864_inl51 && !c866_inl51) && !c868_inl51) && !c870_inl51) && c872_inl51); */
        /* c1088_inl51 <= (((((!c864_inl51 && !c866_inl51) && !c868_inl51) && !c870_inl51) && !c872_inl51) && c874_inl51); */
        /* c1089_inl51 <= ((((((!c864_inl51 && !c866_inl51) && !c868_inl51) && !c870_inl51) && !c872_inl51) && !c874_inl51) && c876_inl51); */
        /* c1090_inl51 <= ((((((!c864_inl51 && !c866_inl51) && !c868_inl51) && !c870_inl51) && !c872_inl51) && !c874_inl51) && !c876_inl51); */
        /* c2334 <= ((c2333 || c2332) && c864_inl51); */
        /* c2335 <= ((c2333 || c2332) && c1084_inl51); */
        /* c2336 <= ((c2333 || c2332) && c1085_inl51); */
        /* c2337 <= ((c2333 || c2332) && c1086_inl51); */
        /* c2338 <= ((c2333 || c2332) && c1087_inl51); */
        /* c2339 <= ((c2333 || c2332) && c1088_inl51); */
        /* c2340 <= ((c2333 || c2332) && c1089_inl51); */
        if (c864_inl51) begin
          array998[4] <= 0;
          /* c2944 <= ((c2943 || c2942) && c864_inl51); */
          retro_main_state <= retro_main_L1_b526_S0;
        end else if (c1084_inl51) begin
          array998[4] <= 0;
          /* c2945 <= ((c2943 || c2942) && c1084_inl51); */
          retro_main_state <= retro_main_L1_b526_S0;
        end else if (c1085_inl51) begin
          array998[4] <= 1;
          /* c2946 <= ((c2943 || c2942) && c1085_inl51); */
          retro_main_state <= retro_main_L1_b526_S0;
        end else if (c1086_inl51) begin
          array998[4] <= 0;
          /* c2947 <= ((c2943 || c2942) && c1086_inl51); */
          retro_main_state <= retro_main_L1_b526_S0;
        end else if (c1087_inl51) begin
          array998[4] <= 0;
          /* c2948 <= ((c2943 || c2942) && c1087_inl51); */
          retro_main_state <= retro_main_L1_b526_S0;
        end else if (c1088_inl51) begin
          array998[4] <= 0;
          /* c2949 <= ((c2943 || c2942) && c1088_inl51); */
          retro_main_state <= retro_main_L1_b526_S0;
        end else if (c1089_inl51) begin
          array998[4] <= 0;
          /* c2950 <= ((c2943 || c2942) && c1089_inl51); */
          retro_main_state <= retro_main_L1_b526_S0;
        end else if (c1090_inl51) begin
          t877_inl51 <= array998[4];
          /* c2951 <= ((c2943 || c2942) && c1090_inl51); */
          /* c2341 <= ((c2333 || c2332) && c1090_inl51); */
          retro_main_state <= retro_main_L1_b526_S1;
        end
      end
      retro_main_L1_b526_S0: begin
        t877_inl51 <= array998[4];
        /* c2951 <= ((c2943 || c2942) && c1090_inl51); */
        /* c2341 <= ((c2333 || c2332) && c1090_inl51); */
        retro_main_state <= retro_main_L1_b526_S1;
      end
      retro_main_L1_b526_S1: begin
        /* c878_inl51 <= (t877_inl51 == -8); */
        /* c2342 <= ((((((((c2341 || c2336) || c2334) || c2335) || c2340) || c2339) || c2338) || c2337) && c878_inl51); */
        if (c878_inl51) begin
          array998[4] <= 0;
          /* c2952 <= ((((((((c2951 || c2946) || c2944) || c2945) || c2950) || c2949) || c2948) || c2947) && c878_inl51); */
          retro_main_state <= retro_main_L1_b528_S0;
        end else begin
          t879_inl51 <= array998[5];
          t881_inl51 <= array998[5];
          t883_inl51 <= array998[5];
          t885_inl51 <= array998[5];
          t887_inl51 <= array998[5];
          t889_inl51 <= array998[5];
          t891_inl51 <= array998[5];
          t893_inl51 <= array998[5];
          t895_inl51 <= array998[5];
          t897_inl51 <= array998[5];
          t899_inl51 <= array998[5];
          t901_inl51 <= array998[5];
          t903_inl51 <= array998[5];
          t905_inl51 <= array998[5];
          t907_inl51 <= array998[5];
          /* c2953 <= ((((((((c2951 || c2946) || c2944) || c2945) || c2950) || c2949) || c2948) || c2947) && !c878_inl51); */
          /* c2343 <= ((((((((c2341 || c2336) || c2334) || c2335) || c2340) || c2339) || c2338) || c2337) && !c878_inl51); */
          retro_main_state <= retro_main_L1_b528_S1;
        end
      end
      retro_main_L1_b528_S0: begin
        t879_inl51 <= array998[5];
        t881_inl51 <= array998[5];
        t883_inl51 <= array998[5];
        t885_inl51 <= array998[5];
        t887_inl51 <= array998[5];
        t889_inl51 <= array998[5];
        t891_inl51 <= array998[5];
        t893_inl51 <= array998[5];
        t895_inl51 <= array998[5];
        t897_inl51 <= array998[5];
        t899_inl51 <= array998[5];
        t901_inl51 <= array998[5];
        t903_inl51 <= array998[5];
        t905_inl51 <= array998[5];
        t907_inl51 <= array998[5];
        /* c2953 <= ((((((((c2951 || c2946) || c2944) || c2945) || c2950) || c2949) || c2948) || c2947) && !c878_inl51); */
        /* c2343 <= ((((((((c2341 || c2336) || c2334) || c2335) || c2340) || c2339) || c2338) || c2337) && !c878_inl51); */
        retro_main_state <= retro_main_L1_b528_S1;
      end
      retro_main_L1_b528_S1: begin
        /* c880_inl51 <= (t879_inl51 == -1); */
        /* c882_inl51 <= (t881_inl51 == -2); */
        /* c884_inl51 <= (t883_inl51 == -3); */
        /* c886_inl51 <= (t885_inl51 == -4); */
        /* c888_inl51 <= (t887_inl51 == -5); */
        /* c890_inl51 <= (t889_inl51 == -6); */
        /* c892_inl51 <= (t891_inl51 == -7); */
        /* c894_inl51 <= (t893_inl51 == -8); */
        /* c896_inl51 <= (t895_inl51 == -9); */
        /* c898_inl51 <= (t897_inl51 == -10); */
        /* c900_inl51 <= (t899_inl51 == -11); */
        /* c902_inl51 <= (t901_inl51 == -12); */
        /* c904_inl51 <= (t903_inl51 == -13); */
        /* c906_inl51 <= (t905_inl51 == -14); */
        /* c908_inl51 <= (t907_inl51 == -15); */
        /* c1091_inl51 <= (!c880_inl51 && c882_inl51); */
        /* c1092_inl51 <= ((!c880_inl51 && !c882_inl51) && c884_inl51); */
        /* c1093_inl51 <= (((!c880_inl51 && !c882_inl51) && !c884_inl51) && c886_inl51); */
        /* c1094_inl51 <= ((((!c880_inl51 && !c882_inl51) && !c884_inl51) && !c886_inl51) && c888_inl51); */
        /* c1095_inl51 <= (((((!c880_inl51 && !c882_inl51) && !c884_inl51) && !c886_inl51) && !c888_inl51) && c890_inl51); */
        /* c1096_inl51 <= ((((((!c880_inl51 && !c882_inl51) && !c884_inl51) && !c886_inl51) && !c888_inl51) && !c890_inl51) && c892_inl51); */
        /* c1097_inl51 <= (((((((!c880_inl51 && !c882_inl51) && !c884_inl51) && !c886_inl51) && !c888_inl51) && !c890_inl51) && !c892_inl51) && c894_inl51); */
        /* c1098_inl51 <= ((((((((!c880_inl51 && !c882_inl51) && !c884_inl51) && !c886_inl51) && !c888_inl51) && !c890_inl51) && !c892_inl51) && !c894_inl51) && c896_inl51); */
        /* c1099_inl51 <= (((((((((!c880_inl51 && !c882_inl51) && !c884_inl51) && !c886_inl51) && !c888_inl51) && !c890_inl51) && !c892_inl51) && !c894_inl51) && !c896_inl51) && c898_inl51); */
        /* c1100_inl51 <= ((((((((((!c880_inl51 && !c882_inl51) && !c884_inl51) && !c886_inl51) && !c888_inl51) && !c890_inl51) && !c892_inl51) && !c894_inl51) && !c896_inl51) && !c898_inl51) && c900_inl51); */
        /* c1101_inl51 <= (((((((((((!c880_inl51 && !c882_inl51) && !c884_inl51) && !c886_inl51) && !c888_inl51) && !c890_inl51) && !c892_inl51) && !c894_inl51) && !c896_inl51) && !c898_inl51) && !c900_inl51) && c902_inl51); */
        /* c1102_inl51 <= ((((((((((((!c880_inl51 && !c882_inl51) && !c884_inl51) && !c886_inl51) && !c888_inl51) && !c890_inl51) && !c892_inl51) && !c894_inl51) && !c896_inl51) && !c898_inl51) && !c900_inl51) && !c902_inl51) && c904_inl51); */
        /* c1103_inl51 <= (((((((((((((!c880_inl51 && !c882_inl51) && !c884_inl51) && !c886_inl51) && !c888_inl51) && !c890_inl51) && !c892_inl51) && !c894_inl51) && !c896_inl51) && !c898_inl51) && !c900_inl51) && !c902_inl51) && !c904_inl51) && c906_inl51); */
        /* c1104_inl51 <= ((((((((((((((!c880_inl51 && !c882_inl51) && !c884_inl51) && !c886_inl51) && !c888_inl51) && !c890_inl51) && !c892_inl51) && !c894_inl51) && !c896_inl51) && !c898_inl51) && !c900_inl51) && !c902_inl51) && !c904_inl51) && !c906_inl51) && c908_inl51); */
        /* c1105_inl51 <= ((((((((((((((!c880_inl51 && !c882_inl51) && !c884_inl51) && !c886_inl51) && !c888_inl51) && !c890_inl51) && !c892_inl51) && !c894_inl51) && !c896_inl51) && !c898_inl51) && !c900_inl51) && !c902_inl51) && !c904_inl51) && !c906_inl51) && !c908_inl51); */
        /* c2344 <= ((c2343 || c2342) && c880_inl51); */
        /* c2345 <= ((c2343 || c2342) && c1091_inl51); */
        /* c2346 <= ((c2343 || c2342) && c1092_inl51); */
        /* c2347 <= ((c2343 || c2342) && c1093_inl51); */
        /* c2348 <= ((c2343 || c2342) && c1094_inl51); */
        /* c2349 <= ((c2343 || c2342) && c1095_inl51); */
        /* c2350 <= ((c2343 || c2342) && c1096_inl51); */
        /* c2351 <= ((c2343 || c2342) && c1097_inl51); */
        /* c2352 <= ((c2343 || c2342) && c1098_inl51); */
        /* c2353 <= ((c2343 || c2342) && c1099_inl51); */
        /* c2354 <= ((c2343 || c2342) && c1100_inl51); */
        /* c2355 <= ((c2343 || c2342) && c1101_inl51); */
        /* c2356 <= ((c2343 || c2342) && c1102_inl51); */
        /* c2357 <= ((c2343 || c2342) && c1103_inl51); */
        /* c2358 <= ((c2343 || c2342) && c1104_inl51); */
        if (c880_inl51) begin
          array998[5] <= 99999;
          /* c2954 <= ((c2953 || c2952) && c880_inl51); */
          retro_main_state <= retro_main_L1_b530_S0;
        end else if (c1091_inl51) begin
          array998[5] <= 0;
          /* c2955 <= ((c2953 || c2952) && c1091_inl51); */
          retro_main_state <= retro_main_L1_b530_S0;
        end else if (c1092_inl51) begin
          array998[5] <= 0;
          /* c2956 <= ((c2953 || c2952) && c1092_inl51); */
          retro_main_state <= retro_main_L1_b530_S0;
        end else if (c1093_inl51) begin
          array998[5] <= 0;
          /* c2957 <= ((c2953 || c2952) && c1093_inl51); */
          retro_main_state <= retro_main_L1_b530_S0;
        end else if (c1094_inl51) begin
          array998[5] <= 128;
          /* c2958 <= ((c2953 || c2952) && c1094_inl51); */
          retro_main_state <= retro_main_L1_b530_S0;
        end else if (c1095_inl51) begin
          array998[5] <= 1024;
          /* c2959 <= ((c2953 || c2952) && c1095_inl51); */
          retro_main_state <= retro_main_L1_b530_S0;
        end else if (c1096_inl51) begin
          array998[5] <= 0;
          /* c2960 <= ((c2953 || c2952) && c1096_inl51); */
          retro_main_state <= retro_main_L1_b530_S0;
        end else if (c1097_inl51) begin
          array998[5] <= 0;
          /* c2961 <= ((c2953 || c2952) && c1097_inl51); */
          retro_main_state <= retro_main_L1_b530_S0;
        end else if (c1098_inl51) begin
          array998[5] <= 0;
          /* c2962 <= ((c2953 || c2952) && c1098_inl51); */
          retro_main_state <= retro_main_L1_b530_S0;
        end else if (c1099_inl51) begin
          array998[5] <= 0;
          /* c2963 <= ((c2953 || c2952) && c1099_inl51); */
          retro_main_state <= retro_main_L1_b530_S0;
        end else if (c1100_inl51) begin
          array998[5] <= 0;
          /* c2964 <= ((c2953 || c2952) && c1100_inl51); */
          retro_main_state <= retro_main_L1_b530_S0;
        end else if (c1101_inl51) begin
          array998[5] <= 0;
          /* c2965 <= ((c2953 || c2952) && c1101_inl51); */
          retro_main_state <= retro_main_L1_b530_S0;
        end else if (c1102_inl51) begin
          array998[5] <= 32;
          /* c2966 <= ((c2953 || c2952) && c1102_inl51); */
          retro_main_state <= retro_main_L1_b530_S0;
        end else if (c1103_inl51) begin
          array998[5] <= 0;
          /* c2967 <= ((c2953 || c2952) && c1103_inl51); */
          retro_main_state <= retro_main_L1_b530_S0;
        end else if (c1104_inl51) begin
          array998[5] <= -1;
          /* c2968 <= ((c2953 || c2952) && c1104_inl51); */
          retro_main_state <= retro_main_L1_b530_S0;
        end else if (c1105_inl51) begin
          t909_inl51 <= array998[8];
          /* c2969 <= ((c2953 || c2952) && c1105_inl51); */
          /* c2359 <= ((c2343 || c2342) && c1105_inl51); */
          /* ip_inl514 <= c2344 ? ip2 : c2345 ? ip2 : c2346 ? ip2 : c2347 ? ip2 : c2348 ? ip2 : c2349 ? ip2 : c2350 ? ip2 : c2351 ? ip2 : c2352 ? 16384 : c2353 ? ip2 : c2354 ? ip2 : c2355 ? ip2 : c2356 ? ip2 : c2357 ? ip2 : c2358 ? ip2 : ((c2343 || c2342) && c1105_inl51) ? ip2 : 'bz; */
          retro_main_state <= retro_main_L1_b530_S1;
        end
      end
      retro_main_L1_b530_S0: begin
        t909_inl51 <= array998[8];
        /* c2969 <= ((c2953 || c2952) && c1105_inl51); */
        /* c2359 <= ((c2343 || c2342) && c1105_inl51); */
        /* ip_inl514 <= c2344 ? ip2 : c2345 ? ip2 : c2346 ? ip2 : c2347 ? ip2 : c2348 ? ip2 : c2349 ? ip2 : c2350 ? ip2 : c2351 ? ip2 : c2352 ? 16384 : c2353 ? ip2 : c2354 ? ip2 : c2355 ? ip2 : c2356 ? ip2 : c2357 ? ip2 : c2358 ? ip2 : ((c2343 || c2342) && c1105_inl51) ? ip2 : 'bz; */
        retro_main_state <= retro_main_L1_b530_S1;
      end
      retro_main_L1_b530_S1: begin
        /* c910_inl51 <= (t909_inl51 == 1); */
        /* c2360 <= ((((((((((((((((c2359 || c2349) || c2344) || c2357) || c2348) || c2347) || c2350) || c2351) || c2356) || c2353) || c2355) || c2358) || c2354) || c2346) || c2352) || c2345) && c910_inl51); */
        if (c910_inl51) begin
          array998[8] <= 0;
          /* c2970 <= ((((((((((((((((c2969 || c2959) || c2954) || c2967) || c2958) || c2957) || c2960) || c2961) || c2966) || c2963) || c2965) || c2968) || c2964) || c2956) || c2962) || c2955) && c910_inl51); */
          retro_main_state <= retro_main_L1_b532_S0;
        end else begin
          /* c2971 <= ((((((((((((((((c2969 || c2959) || c2954) || c2967) || c2958) || c2957) || c2960) || c2961) || c2966) || c2963) || c2965) || c2968) || c2964) || c2956) || c2962) || c2955) && !c910_inl51); */
          /* c2361 <= ((((((((((((((((c2359 || c2349) || c2344) || c2357) || c2348) || c2347) || c2350) || c2351) || c2356) || c2353) || c2355) || c2358) || c2354) || c2346) || c2352) || c2345) && !c910_inl51); */
          retro_main_state <= retro_main_L1_b198_S0;
        end
      end
      retro_main_L1_b532_S0: begin
        /* c2971 <= ((((((((((((((((c2969 || c2959) || c2954) || c2967) || c2958) || c2957) || c2960) || c2961) || c2966) || c2963) || c2965) || c2968) || c2964) || c2956) || c2962) || c2955) && !c910_inl51); */
        /* c2361 <= ((((((((((((((((c2359 || c2349) || c2344) || c2357) || c2348) || c2347) || c2350) || c2351) || c2356) || c2353) || c2355) || c2358) || c2354) || c2346) || c2352) || c2345) && !c910_inl51); */
        retro_main_state <= retro_main_L1_b198_S0;
      end
      retro_main_L1_b198_S0: begin
        a6 <= (c2157 && c916) ? a6 : c2159 ? a6 : c2160 ? a6 : c2161 ? a6 : c2162 ? a6 : c2163 ? a6 : c2164 ? a6 : c2246 ? a6 : c2247 ? a6 : c2166 ? a6 : c2167 ? a6 : c2168 ? stack0_top2 : c2169 ? stack0_top2 : c2170 ? stack0_top2 : c2171 ? stack0_top2 : c2172 ? a6 : c2173 ? a6 : c2174 ? a6 : c2175 ? a6 : c2176 ? a6 : (c2286 || c2284) ? a6 : c2178 ? a6 : c2179 ? a6 : c2180 ? a6 : c2181 ? a6 : c2182 ? a6 : c2212 ? a6 : (c2183 && !c964) ? a6 : c2184 ? a6 : c2185 ? a6 : c2186 ? a6 : c2187 ? a6 : (c2361 || c2360) ? a6 : (c2188 && !c967) ? a6 : (c2157 && c1136) ? a6 : c2158 ? a6 : 'bz;
        /* address0_pos8 <= (c2157 && c916) ? address0_pos2 : c2159 ? address0_pos2 : c2160 ? address0_pos2 : c2161 ? address0_pos2 : c2162 ? address0_pos2 : c2163 ? address0_pos3 : c2164 ? address0_pos4 : c2246 ? address0_pos2 : c2247 ? address0_pos2 : c2166 ? address0_pos2 : c2167 ? address0_pos5 : c2168 ? address0_pos2 : c2169 ? address0_pos2 : c2170 ? address0_pos2 : c2171 ? address0_pos2 : c2172 ? address0_pos2 : c2173 ? address0_pos2 : c2174 ? address0_pos2 : c2175 ? address0_pos2 : c2176 ? address0_pos2 : (c2286 || c2284) ? address0_pos2 : c2178 ? address0_pos2 : c2179 ? address0_pos2 : c2180 ? address0_pos2 : c2181 ? address0_pos2 : c2182 ? address0_pos2 : c2212 ? address0_pos6 : (c2183 && !c964) ? address0_pos2 : c2184 ? address0_pos2 : c2185 ? address0_pos2 : c2186 ? address0_pos2 : c2187 ? address0_pos2 : (c2361 || c2360) ? address0_pos2 : (c2188 && !c967) ? address0_pos2 : (c2157 && c1136) ? address0_pos2 : c2158 ? address0_pos7 : 'bz; */
        /* address0_second8 <= (c2157 && c916) ? address0_second2 : c2159 ? address0_second2 : c2160 ? address0_second2 : c2161 ? address0_second2 : c2162 ? address0_second2 : c2163 ? address0_top2 : c2164 ? address0_second4 : c2246 ? address0_second2 : c2247 ? address0_second2 : c2166 ? address0_second2 : c2167 ? address0_second5 : c2168 ? address0_second2 : c2169 ? address0_second2 : c2170 ? address0_second2 : c2171 ? address0_second2 : c2172 ? address0_second2 : c2173 ? address0_second2 : c2174 ? address0_second2 : c2175 ? address0_second2 : c2176 ? address0_second2 : (c2286 || c2284) ? address0_second2 : c2178 ? address0_second2 : c2179 ? address0_second2 : c2180 ? address0_second2 : c2181 ? address0_second2 : c2182 ? address0_second2 : c2212 ? address0_second6 : (c2183 && !c964) ? address0_second2 : c2184 ? address0_second2 : c2185 ? address0_second2 : c2186 ? address0_second2 : c2187 ? address0_second2 : (c2361 || c2360) ? address0_second2 : (c2188 && !c967) ? address0_second2 : (c2157 && c1136) ? address0_second2 : c2158 ? address0_top2 : 'bz; */
        /* address0_top8 <= (c2157 && c916) ? address0_top2 : c2159 ? address0_top2 : c2160 ? address0_top2 : c2161 ? address0_top2 : c2162 ? address0_top2 : c2163 ? stack0_top2 : c2164 ? address0_second2 : c2246 ? address0_top2 : c2247 ? address0_top2 : c2166 ? address0_top2 : c2167 ? address0_second2 : c2168 ? address0_top2 : c2169 ? address0_top2 : c2170 ? address0_top2 : c2171 ? address0_top2 : c2172 ? address0_top2 : c2173 ? address0_top2 : c2174 ? address0_top2 : c2175 ? address0_top2 : c2176 ? address0_top2 : (c2286 || c2284) ? address0_top2 : c2178 ? address0_top2 : c2179 ? address0_top2 : c2180 ? address0_top2 : c2181 ? address0_top2 : c2182 ? address0_top2 : c2212 ? address0_second2 : (c2183 && !c964) ? address0_top2 : c2184 ? address0_top2 : c2185 ? address0_top2 : c2186 ? address0_top2 : c2187 ? address0_top2 : (c2361 || c2360) ? address0_top2 : (c2188 && !c967) ? address0_top2 : (c2157 && c1136) ? address0_top2 : c2158 ? ip2 : 'bz; */
        b6 <= (c2157 && c916) ? b6 : c2159 ? b6 : c2160 ? b6 : c2161 ? b6 : c2162 ? b6 : c2163 ? b6 : c2164 ? b6 : c2246 ? b6 : c2247 ? b6 : c2166 ? b6 : c2167 ? b6 : c2168 ? stack0_second2 : c2169 ? stack0_second2 : c2170 ? stack0_second2 : c2171 ? stack0_second2 : c2172 ? b6 : c2173 ? b6 : c2174 ? b6 : c2175 ? b6 : c2176 ? b6 : (c2286 || c2284) ? b6 : c2178 ? b6 : c2179 ? b6 : c2180 ? b6 : c2181 ? b6 : c2182 ? b6 : c2212 ? b6 : (c2183 && !c964) ? b6 : c2184 ? b6 : c2185 ? b6 : c2186 ? b6 : c2187 ? b6 : (c2361 || c2360) ? b6 : (c2188 && !c967) ? b6 : (c2157 && c1136) ? b6 : c2158 ? b6 : 'bz;
        /* ip21 <= (c2157 && c916) ? ip2 : c2159 ? ip3 : c2160 ? ip2 : c2161 ? ip2 : c2162 ? ip2 : c2163 ? ip2 : c2164 ? ip2 : c2246 ? ip5 : c2247 ? ip6 : c2166 ? ip8 : c2167 ? address0_top2 : c2168 ? t2660 : c2169 ? t2670 : c2170 ? t2680 : c2171 ? t2690 : c2172 ? ip2 : c2173 ? ip2 : c2174 ? ip2 : c2175 ? ip2 : c2176 ? ip2 : (c2286 || c2284) ? ip2 : c2178 ? ip2 : c2179 ? ip2 : c2180 ? ip2 : c2181 ? ip2 : c2182 ? ip2 : c2212 ? address0_top2 : (c2183 && !c964) ? ip2 : c2184 ? ip2 : c2185 ? ip2 : c2186 ? ip2 : c2187 ? ip2 : (c2361 || c2360) ? ip_inl514 : (c2188 && !c967) ? ip2 : (c2157 && c1136) ? ip2 : c2158 ? ip20 : 'bz; */
        /* stack0_pos35 <= (c2157 && c916) ? stack0_pos2 : c2159 ? stack0_pos3 : c2160 ? stack0_pos4 : c2161 ? stack0_pos5 : c2162 ? stack0_pos2 : c2163 ? stack0_pos6 : c2164 ? stack0_pos7 : c2246 ? stack0_pos2 : c2247 ? stack0_pos8 : c2166 ? stack0_pos2 : c2167 ? stack0_pos2 : c2168 ? stack0_pos10 : c2169 ? stack0_pos12 : c2170 ? stack0_pos14 : c2171 ? stack0_pos16 : c2172 ? stack0_pos2 : c2173 ? stack0_pos18 : c2174 ? stack0_pos19 : c2175 ? stack0_pos20 : c2176 ? stack0_pos21 : (c2286 || c2284) ? stack0_pos2 : c2178 ? stack0_pos22 : c2179 ? stack0_pos23 : c2180 ? stack0_pos24 : c2181 ? stack0_pos25 : c2182 ? stack0_pos26 : c2212 ? stack0_pos27 : (c2183 && !c964) ? stack0_pos2 : c2184 ? stack0_pos2 : c2185 ? stack0_pos2 : c2186 ? stack0_pos2 : c2187 ? stack0_pos29 : (c2361 || c2360) ? stack0_pos34 : (c2188 && !c967) ? stack0_pos2 : (c2157 && c1136) ? stack0_pos2 : c2158 ? stack0_pos2 : 'bz; */
        /* stack0_second37 <= (c2157 && c916) ? stack0_second2 : c2159 ? stack0_top2 : c2160 ? stack0_top2 : c2161 ? stack0_second5 : c2162 ? stack0_top2 : c2163 ? stack0_second7 : c2164 ? stack0_top2 : c2246 ? stack0_second2 : c2247 ? stack0_second9 : c2166 ? stack0_second2 : c2167 ? stack0_second2 : c2168 ? stack0_second11 : c2169 ? stack0_second13 : c2170 ? stack0_second15 : c2171 ? stack0_second17 : c2172 ? stack0_second2 : c2173 ? stack0_second19 : c2174 ? stack0_second20 : c2175 ? stack0_second21 : c2176 ? stack0_second22 : (c2286 || c2284) ? stack0_second23 : c2178 ? stack0_second24 : c2179 ? stack0_second25 : c2180 ? stack0_second26 : c2181 ? stack0_second27 : c2182 ? stack0_second28 : c2212 ? stack0_second29 : (c2183 && !c964) ? stack0_second2 : c2184 ? stack0_second2 : c2185 ? stack0_second2 : c2186 ? stack0_second2 : c2187 ? stack0_second31 : (c2361 || c2360) ? stack0_second36 : (c2188 && !c967) ? stack0_second2 : (c2157 && c1136) ? stack0_second2 : c2158 ? stack0_second2 : 'bz; */
        /* stack0_top50 <= (c2157 && c916) ? stack0_top2 : c2159 ? t947 : c2160 ? stack0_top2 : c2161 ? stack0_second2 : c2162 ? stack0_second2 : c2163 ? stack0_second2 : c2164 ? address0_top2 : c2246 ? stack0_top9 : c2247 ? stack0_second2 : c2166 ? stack0_top2 : c2167 ? stack0_top2 : c2168 ? stack0_second10 : c2169 ? stack0_second12 : c2170 ? stack0_second14 : c2171 ? stack0_second16 : c2172 ? stack0_top19 : c2173 ? stack0_second18 : c2174 ? stack0_top23 : c2175 ? stack0_top25 : c2176 ? stack0_top27 : (c2286 || c2284) ? stack0_top28 : c2178 ? stack0_top30 : c2179 ? stack0_top32 : c2180 ? stack0_top34 : c2181 ? stack0_top36 : c2182 ? stack0_top38 : c2212 ? stack0_second2 : (c2183 && !c964) ? stack0_top2 : c2184 ? stack0_top40 : c2185 ? stack0_top41 : c2186 ? stack0_top42 : c2187 ? stack0_second30 : (c2361 || c2360) ? stack0_top49 : (c2188 && !c967) ? stack0_top2 : (c2157 && c1136) ? stack0_top2 : c2158 ? stack0_top2 : 'bz; */
        t11 <= (c2157 && c916) ? t11 : c2159 ? t11 : c2160 ? t11 : c2161 ? t11 : c2162 ? t11 : c2163 ? t11 : c2164 ? t11 : c2246 ? t11 : c2247 ? t11 : c2166 ? t11 : c2167 ? t11 : c2168 ? t11 : c2169 ? t11 : c2170 ? t11 : c2171 ? t11 : c2172 ? t11 : c2173 ? t11 : c2174 ? stack0_top2 : c2175 ? stack0_top2 : c2176 ? stack0_top2 : (c2286 || c2284) ? t11 : c2178 ? stack0_top2 : c2179 ? stack0_top2 : c2180 ? stack0_top2 : c2181 ? stack0_top2 : c2182 ? stack0_top2 : c2212 ? t11 : (c2183 && !c964) ? t11 : c2184 ? t11 : c2185 ? t11 : c2186 ? stack0_top2 : c2187 ? t11 : (c2361 || c2360) ? t11 : (c2188 && !c967) ? t11 : (c2157 && c1136) ? t11 : c2158 ? t11 : 'bz;
        /* ip22 <= (ip21 + 1); */
        address0_pos2 <= address0_pos8;
        address0_second2 <= address0_second8;
        stack0_pos2 <= stack0_pos35;
        stack0_second2 <= stack0_second37;
        address0_top2 <= address0_top8;
        ip2 <= ip22;
        stack0_top2 <= stack0_top50;
        retro_main_state <= retro_main_L1_b198_S1;
      end
      retro_main_L1_b198_S1: begin
        retro_main_state <= retro_main_L1_while2_S0;
      end
      retro_main_L10_while463_S0: begin
        io_ports_addr <= 1;
        io_ports_we <= 0;
        io_ports_req <= 1;
        retro_main_state <= retro_main_L10_while463_S1;
      end
      retro_main_L10_while463_S1: begin
        /*wait for output of io_ports*/
        retro_main_state <= retro_main_L10_while463_S2;
      end
      retro_main_L10_while463_S2: begin
        t983_inl3_inl5_inl51 <= io_ports_q;
        io_ports_req <= 0;
        retro_main_state <= retro_main_L10_while463_S3;
      end
      retro_main_L10_while463_S3: begin
        /* cmd_reply_inl3_inl5_inl51 <= (t983_inl3_inl5_inl51 & 4294967295); */
        /* c985_inl3_inl5_inl51 <= (cmd_reply_inl3_inl5_inl51 == 2147483648); */
        if (c985_inl3_inl5_inl51) begin
          io_ports_addr <= 0;
          io_ports_we <= 0;
          io_ports_req <= 1;
          retro_main_state <= retro_main_L11_while470_S1;
        end else begin
          /* c2925 <= (c2919 && !c985_inl3_inl5_inl51); */
          /* c2314 <= (c2300 && !c985_inl3_inl5_inl51); */
          retro_main_state <= retro_main_L10_while463_S0;
        end
      end
      retro_main_L11_while470_S0: begin
        io_ports_addr <= 0;
        io_ports_we <= 0;
        io_ports_req <= 1;
        retro_main_state <= retro_main_L11_while470_S1;
      end
      retro_main_L11_while470_S1: begin
        /*wait for output of io_ports*/
        retro_main_state <= retro_main_L11_while470_S2;
      end
      retro_main_L11_while470_S2: begin
        t992_inl1_inl6_inl51 <= io_ports_q;
        io_ports_req <= 0;
        retro_main_state <= retro_main_L11_while470_S3;
      end
      retro_main_L11_while470_S3: begin
        /* cmd_reply_inl1_inl6_inl51 <= (t992_inl1_inl6_inl51 & 4294967295); */
        /* t993_inl1_inl6_inl51 <= (cmd_reply_inl1_inl6_inl51 & 2147483648); */
        /* c994_inl1_inl6_inl51 <= (t993_inl1_inl6_inl51 == 0); */
        if (c994_inl1_inl6_inl51) begin
          io_ports_addr <= 3;
          io_ports_we <= 1;
          io_ports_req <= 1;
          io_ports_d <= 32;
          retro_main_state <= retro_main_L1_whileexit472_S1;
        end else begin
          /* c2927 <= (c2919 && !c994_inl1_inl6_inl51); */
          /* c2316 <= (c2300 && !c994_inl1_inl6_inl51); */
          retro_main_state <= retro_main_L11_while470_S0;
        end
      end
      retro_main_L12_while475_S0: begin
        io_ports_addr <= 1;
        io_ports_we <= 0;
        io_ports_req <= 1;
        retro_main_state <= retro_main_L12_while475_S1;
      end
      retro_main_L12_while475_S1: begin
        /*wait for output of io_ports*/
        retro_main_state <= retro_main_L12_while475_S2;
      end
      retro_main_L12_while475_S2: begin
        t983_inl2_inl6_inl51 <= io_ports_q;
        io_ports_req <= 0;
        retro_main_state <= retro_main_L12_while475_S3;
      end
      retro_main_L12_while475_S3: begin
        /* cmd_reply_inl2_inl6_inl51 <= (t983_inl2_inl6_inl51 & 4294967295); */
        /* c985_inl2_inl6_inl51 <= (cmd_reply_inl2_inl6_inl51 == 2147483649); */
        if (c985_inl2_inl6_inl51) begin
          io_ports_addr <= 1;
          io_ports_we <= 1;
          io_ports_req <= 1;
          io_ports_d <= 0;
          retro_main_state <= retro_main_L1_whileexit477_S1;
        end else begin
          /* c2928 <= (c2919 && !c985_inl2_inl6_inl51); */
          /* c2317 <= (c2300 && !c985_inl2_inl6_inl51); */
          retro_main_state <= retro_main_L12_while475_S0;
        end
      end
      retro_main_L13_while480_S0: begin
        io_ports_addr <= 1;
        io_ports_we <= 0;
        io_ports_req <= 1;
        retro_main_state <= retro_main_L13_while480_S1;
      end
      retro_main_L13_while480_S1: begin
        /*wait for output of io_ports*/
        retro_main_state <= retro_main_L13_while480_S2;
      end
      retro_main_L13_while480_S2: begin
        t983_inl3_inl6_inl51 <= io_ports_q;
        io_ports_req <= 0;
        retro_main_state <= retro_main_L13_while480_S3;
      end
      retro_main_L13_while480_S3: begin
        /* cmd_reply_inl3_inl6_inl51 <= (t983_inl3_inl6_inl51 & 4294967295); */
        /* c985_inl3_inl6_inl51 <= (cmd_reply_inl3_inl6_inl51 == 2147483648); */
        if (c985_inl3_inl6_inl51) begin
          io_ports_addr <= 0;
          io_ports_we <= 0;
          io_ports_req <= 1;
          retro_main_state <= retro_main_L14_while487_S1;
        end else begin
          /* c2929 <= (c2919 && !c985_inl3_inl6_inl51); */
          /* c2318 <= (c2300 && !c985_inl3_inl6_inl51); */
          retro_main_state <= retro_main_L13_while480_S0;
        end
      end
      retro_main_L14_while487_S0: begin
        io_ports_addr <= 0;
        io_ports_we <= 0;
        io_ports_req <= 1;
        retro_main_state <= retro_main_L14_while487_S1;
      end
      retro_main_L14_while487_S1: begin
        /*wait for output of io_ports*/
        retro_main_state <= retro_main_L14_while487_S2;
      end
      retro_main_L14_while487_S2: begin
        t992_inl1_inl7_inl51 <= io_ports_q;
        io_ports_req <= 0;
        retro_main_state <= retro_main_L14_while487_S3;
      end
      retro_main_L14_while487_S3: begin
        /* cmd_reply_inl1_inl7_inl51 <= (t992_inl1_inl7_inl51 & 4294967295); */
        /* t993_inl1_inl7_inl51 <= (cmd_reply_inl1_inl7_inl51 & 2147483648); */
        /* c994_inl1_inl7_inl51 <= (t993_inl1_inl7_inl51 == 0); */
        if (c994_inl1_inl7_inl51) begin
          io_ports_addr <= 3;
          io_ports_we <= 1;
          io_ports_req <= 1;
          io_ports_d <= 8;
          retro_main_state <= retro_main_L1_whileexit489_S1;
        end else begin
          /* c2930 <= (c2919 && !c994_inl1_inl7_inl51); */
          /* c2319 <= (c2300 && !c994_inl1_inl7_inl51); */
          retro_main_state <= retro_main_L14_while487_S0;
        end
      end
      retro_main_L15_while492_S0: begin
        io_ports_addr <= 1;
        io_ports_we <= 0;
        io_ports_req <= 1;
        retro_main_state <= retro_main_L15_while492_S1;
      end
      retro_main_L15_while492_S1: begin
        /*wait for output of io_ports*/
        retro_main_state <= retro_main_L15_while492_S2;
      end
      retro_main_L15_while492_S2: begin
        t983_inl2_inl7_inl51 <= io_ports_q;
        io_ports_req <= 0;
        retro_main_state <= retro_main_L15_while492_S3;
      end
      retro_main_L15_while492_S3: begin
        /* cmd_reply_inl2_inl7_inl51 <= (t983_inl2_inl7_inl51 & 4294967295); */
        /* c985_inl2_inl7_inl51 <= (cmd_reply_inl2_inl7_inl51 == 2147483649); */
        if (c985_inl2_inl7_inl51) begin
          io_ports_addr <= 1;
          io_ports_we <= 1;
          io_ports_req <= 1;
          io_ports_d <= 0;
          retro_main_state <= retro_main_L1_whileexit494_S1;
        end else begin
          /* c2931 <= (c2919 && !c985_inl2_inl7_inl51); */
          /* c2320 <= (c2300 && !c985_inl2_inl7_inl51); */
          retro_main_state <= retro_main_L15_while492_S0;
        end
      end
      retro_main_L16_while497_S0: begin
        io_ports_addr <= 1;
        io_ports_we <= 0;
        io_ports_req <= 1;
        retro_main_state <= retro_main_L16_while497_S1;
      end
      retro_main_L16_while497_S1: begin
        /*wait for output of io_ports*/
        retro_main_state <= retro_main_L16_while497_S2;
      end
      retro_main_L16_while497_S2: begin
        t983_inl3_inl7_inl51 <= io_ports_q;
        io_ports_req <= 0;
        retro_main_state <= retro_main_L16_while497_S3;
      end
      retro_main_L16_while497_S3: begin
        /* cmd_reply_inl3_inl7_inl51 <= (t983_inl3_inl7_inl51 & 4294967295); */
        /* c985_inl3_inl7_inl51 <= (cmd_reply_inl3_inl7_inl51 == 2147483648); */
        if (c985_inl3_inl7_inl51) begin
          /* stack0_pos33 <= (c2300 && c985_inl3_inl7_inl51) ? stack0_pos30 : (c2301 && c985_inl3_inl8_inl51) ? stack0_pos31 : c2298 ? stack0_pos32 : 'bz; */
          /* c2932 <= (c2920 && c985_inl3_inl8_inl51); */
          /* c2933 <= (c2919 && c985_inl3_inl7_inl51); */
          /* stack0_second35 <= (c2300 && c985_inl3_inl7_inl51) ? stack0_second32 : (c2301 && c985_inl3_inl8_inl51) ? stack0_second33 : c2298 ? stack0_second34 : 'bz; */
          /* c2322 <= (c2301 && c985_inl3_inl8_inl51); */
          /* c2323 <= (c2300 && c985_inl3_inl7_inl51); */
          retro_main_state <= retro_main_L17_while505_S0;
        end else begin
          /* c2934 <= (c2919 && !c985_inl3_inl7_inl51); */
          /* c2324 <= (c2300 && !c985_inl3_inl7_inl51); */
          retro_main_state <= retro_main_L16_while497_S0;
        end
      end
      retro_main_L17_while505_S0: begin
        io_ports_addr <= 0;
        io_ports_we <= 0;
        io_ports_req <= 1;
        retro_main_state <= retro_main_L17_while505_S1;
      end
      retro_main_L17_while505_S1: begin
        /*wait for output of io_ports*/
        retro_main_state <= retro_main_L17_while505_S2;
      end
      retro_main_L17_while505_S2: begin
        t992_inl1_inl9_inl51 <= io_ports_q;
        io_ports_req <= 0;
        retro_main_state <= retro_main_L17_while505_S3;
      end
      retro_main_L17_while505_S3: begin
        /* cmd_reply_inl1_inl9_inl51 <= (t992_inl1_inl9_inl51 & 4294967295); */
        /* t993_inl1_inl9_inl51 <= (cmd_reply_inl1_inl9_inl51 & 2147483648); */
        /* c994_inl1_inl9_inl51 <= (t993_inl1_inl9_inl51 == 0); */
        if (c994_inl1_inl9_inl51) begin
          io_ports_addr <= 1;
          io_ports_we <= 1;
          io_ports_req <= 1;
          io_ports_d <= 3;
          retro_main_state <= retro_main_L1_whileexit507_S1;
        end else begin
          /* c2935 <= (((c2918 || c2932) || c2933) && !c994_inl1_inl9_inl51); */
          /* c2325 <= (((c2298 || c2322) || c2323) && !c994_inl1_inl9_inl51); */
          retro_main_state <= retro_main_L17_while505_S0;
        end
      end
      retro_main_L18_while510_S0: begin
        io_ports_addr <= 1;
        io_ports_we <= 0;
        io_ports_req <= 1;
        retro_main_state <= retro_main_L18_while510_S1;
      end
      retro_main_L18_while510_S1: begin
        /*wait for output of io_ports*/
        retro_main_state <= retro_main_L18_while510_S2;
      end
      retro_main_L18_while510_S2: begin
        t983_inl2_inl9_inl51 <= io_ports_q;
        io_ports_req <= 0;
        retro_main_state <= retro_main_L18_while510_S3;
      end
      retro_main_L18_while510_S3: begin
        /* cmd_reply_inl2_inl9_inl51 <= (t983_inl2_inl9_inl51 & 4294967295); */
        /* c985_inl2_inl9_inl51 <= (cmd_reply_inl2_inl9_inl51 == 2147483651); */
        if (c985_inl2_inl9_inl51) begin
          io_ports_addr <= 1;
          io_ports_we <= 1;
          io_ports_req <= 1;
          io_ports_d <= 0;
          retro_main_state <= retro_main_L1_whileexit512_S1;
        end else begin
          /* c2936 <= (((c2918 || c2932) || c2933) && !c985_inl2_inl9_inl51); */
          /* c2326 <= (((c2298 || c2322) || c2323) && !c985_inl2_inl9_inl51); */
          retro_main_state <= retro_main_L18_while510_S0;
        end
      end
      retro_main_L19_while515_S0: begin
        io_ports_addr <= 1;
        io_ports_we <= 0;
        io_ports_req <= 1;
        retro_main_state <= retro_main_L19_while515_S1;
      end
      retro_main_L19_while515_S1: begin
        /*wait for output of io_ports*/
        retro_main_state <= retro_main_L19_while515_S2;
      end
      retro_main_L19_while515_S2: begin
        t983_inl3_inl9_inl51 <= io_ports_q;
        io_ports_req <= 0;
        retro_main_state <= retro_main_L19_while515_S3;
      end
      retro_main_L19_while515_S3: begin
        /* cmd_reply_inl3_inl9_inl51 <= (t983_inl3_inl9_inl51 & 4294967295); */
        /* c985_inl3_inl9_inl51 <= (cmd_reply_inl3_inl9_inl51 == 2147483648); */
        if (c985_inl3_inl9_inl51) begin
          array998[2] <= 0;
          retro_main_state <= retro_main_L1_b520_S0;
        end else begin
          /* c2937 <= (((c2918 || c2932) || c2933) && !c985_inl3_inl9_inl51); */
          /* c2327 <= (((c2298 || c2322) || c2323) && !c985_inl3_inl9_inl51); */
          retro_main_state <= retro_main_L19_while515_S0;
        end
      end
      retro_main_L2_while427_S0: begin
        io_ports_addr <= 0;
        io_ports_we <= 0;
        io_ports_req <= 1;
        retro_main_state <= retro_main_L2_while427_S1;
      end
      retro_main_L2_while427_S1: begin
        /*wait for output of io_ports*/
        retro_main_state <= retro_main_L2_while427_S2;
      end
      retro_main_L2_while427_S2: begin
        t992_inl1_inl1_inl51 <= io_ports_q;
        io_ports_req <= 0;
        retro_main_state <= retro_main_L2_while427_S3;
      end
      retro_main_L2_while427_S3: begin
        /* cmd_reply_inl1_inl1_inl51 <= (t992_inl1_inl1_inl51 & 4294967295); */
        /* t993_inl1_inl1_inl51 <= (cmd_reply_inl1_inl1_inl51 & 2147483648); */
        /* c994_inl1_inl1_inl51 <= (t993_inl1_inl1_inl51 == 0); */
        if (c994_inl1_inl1_inl51) begin
          io_ports_addr <= 1;
          io_ports_we <= 1;
          io_ports_req <= 1;
          io_ports_d <= 2;
          retro_main_state <= retro_main_L1_whileexit429_S1;
        end else begin
          /* c2905 <= (c2901 && !c994_inl1_inl1_inl51); */
          /* c2275 <= (c2243 && !c994_inl1_inl1_inl51); */
          retro_main_state <= retro_main_L2_while427_S0;
        end
      end
      retro_main_L20_fortest393_S0: begin
        /* c986_inl1_inl49 <= (i_inl1_inl493 < 31); */
        if (c986_inl1_inl49) begin
          /* t987_inl1_inl49 <= (test_bit_inl1_inl493 & x_inl1_inl49); */
          /* c2900 <= (c2876 && c986_inl1_inl49); */
          /* c2235 <= (c2177 && c986_inl1_inl49); */
          /* c988_inl1_inl49 <= (t987_inl1_inl49 != 0); */
          if (c988_inl1_inl49) begin
            /* c2902 <= (c2900 && c988_inl1_inl49); */
            /* c2256 <= (c2235 && c988_inl1_inl49); */
            retro_main_state <= retro_main_L1_exit396_S0;
          end else begin
            /* test_bit_inl1_inl494 <= (test_bit_inl1_inl493 >>> 1); */
            /* n_inl1_inl494 <= (n_inl1_inl493 + 1); */
            /* i_inl1_inl494 <= (i_inl1_inl493 + 1); */
            i_inl1_inl493 <= i_inl1_inl494;
            n_inl1_inl493 <= n_inl1_inl494;
            test_bit_inl1_inl493 <= test_bit_inl1_inl494;
            /* c2903 <= (c2900 && !c988_inl1_inl49); */
            /* c2257 <= (c2235 && !c988_inl1_inl49); */
            retro_main_state <= retro_main_L20_fortest393_S0;
          end
        end else begin
          i_inl2_inl493 <= 0;
          n_inl2_inl493 <= 0;
          test_bit_inl2_inl493 <= 1073741824;
          /* x_inl2_inl49 <= abs_b_inl492; */
          /* c2904 <= (c2876 && !c986_inl1_inl49); */
          retro_main_state <= retro_main_L1_exit396_S1;
        end
      end
      retro_main_L21_fortest399_S0: begin
        /* c986_inl2_inl49 <= (i_inl2_inl493 < 31); */
        if (c986_inl2_inl49) begin
          /* t987_inl2_inl49 <= (test_bit_inl2_inl493 & x_inl2_inl49); */
          /* c2906 <= ((c2904 || c2902) && c986_inl2_inl49); */
          /* c2282 <= ((c2177 || c2256) && c986_inl2_inl49); */
          /* c988_inl2_inl49 <= (t987_inl2_inl49 != 0); */
          if (c988_inl2_inl49) begin
            /* c2908 <= (c2906 && c988_inl2_inl49); */
            /* c2284 <= (c2282 && c988_inl2_inl49); */
            retro_main_state <= retro_main_L1_exit402_S0;
          end else begin
            /* test_bit_inl2_inl494 <= (test_bit_inl2_inl493 >>> 1); */
            /* n_inl2_inl494 <= (n_inl2_inl493 + 1); */
            /* i_inl2_inl494 <= (i_inl2_inl493 + 1); */
            i_inl2_inl493 <= i_inl2_inl494;
            n_inl2_inl493 <= n_inl2_inl494;
            test_bit_inl2_inl493 <= test_bit_inl2_inl494;
            /* c2909 <= (c2906 && !c988_inl2_inl49); */
            /* c2285 <= (c2282 && !c988_inl2_inl49); */
            retro_main_state <= retro_main_L21_fortest399_S0;
          end
        end else begin
          c_bit_inl493 <= 0;
          i_inl493 <= 0;
          abs_a_inl493 <= abs_a_inl492;
          /* find_zero_len_result2_inl494 <= c2284 ? n_inl2_inl493 : (c2177 || c2256) ? 0 : 'bz; */
          /* c2286 <= (c2177 || c2256); */
          /* c2910 <= ((c2904 || c2902) && !c986_inl2_inl49); */
          /* abs_b_inl493 <= (abs_b_inl492 << find_zero_len_result2_inl494); */
          /* t486_inl49 <= (find_zero_len_result2_inl494 + 1); */
          abs_b_inl494 <= abs_b_inl493;
          retro_main_state <= retro_main_L1_exit402_S1;
        end
      end
      retro_main_L22_fortest404_S0: begin
        /* c973_inl49 <= (i_inl493 < t486_inl49); */
        if (c973_inl49) begin
          /* c974_inl49 <= (abs_a_inl493 >= abs_b_inl494); */
          /* c_bit_inl496 <= (c_bit_inl493 << 1); */
          /* abs_a_inl496 <= (abs_a_inl493 - abs_b_inl494); */
          /* c_bit_inl498 <= (c_bit_inl493 << 1); */
          /* abs_b_inl495 <= (abs_b_inl494 >>> 1); */
          /* i_inl494 <= (i_inl493 + 1); */
          /* c2913 <= ((c2910 || c2908) && c973_inl49); */
          /* c2289 <= ((c2286 || c2284) && c973_inl49); */
          /* c_bit_inl497 <= (c_bit_inl496 | 1); */
          i_inl493 <= i_inl494;
          /* c2292 <= (c2289 && c974_inl49); */
          /* c2293 <= (c2289 && !c974_inl49); */
          /* abs_a_inl497 <= c2292 ? abs_a_inl496 : c2293 ? abs_a_inl493 : 'bz; */
          /* c_bit_inl499 <= c2292 ? c_bit_inl497 : c2293 ? c_bit_inl498 : 'bz; */
          abs_a_inl493 <= abs_a_inl497;
          c_bit_inl493 <= c_bit_inl499;
          abs_b_inl494 <= abs_b_inl495;
          retro_main_state <= retro_main_L22_fortest404_S0;
        end else begin
          /* c_bit_inl494 <= (c_bit_inl493 | 2147483648); */
          /* c975_inl49 <= (t970_inl49 != 0); */
          /* abs_a_inl494 <= (abs_a_inl493 | 2147483648); */
          /* t976_inl49 <= (t970_inl49 ^ t972_inl49); */
          /* c977_inl49 <= (t976_inl49 != 0); */
          /* c2294 <= ((c2286 || c2284) && c975_inl49); */
          /* c2296 <= ((c2286 || c2284) && !c975_inl49); */
          /* abs_a_inl495 <= c2294 ? abs_a_inl494 : ((c2286 || c2284) && !c975_inl49) ? abs_a_inl493 : 'bz; */
          /* c2299 <= ((c2296 || c2294) && c977_inl49); */
          /* c_bit_inl495 <= c2299 ? c_bit_inl494 : ((c2296 || c2294) && !c977_inl49) ? c_bit_inl493 : 'bz; */
          array995_inl49[0] <= c_bit_inl495;
          array995_inl49[1] <= abs_a_inl495;
          retro_main_state <= retro_main_L1_forelse409_S2;
        end
      end
      retro_main_L3_while432_S0: begin
        io_ports_addr <= 1;
        io_ports_we <= 0;
        io_ports_req <= 1;
        retro_main_state <= retro_main_L3_while432_S1;
      end
      retro_main_L3_while432_S1: begin
        /*wait for output of io_ports*/
        retro_main_state <= retro_main_L3_while432_S2;
      end
      retro_main_L3_while432_S2: begin
        t983_inl2_inl1_inl51 <= io_ports_q;
        io_ports_req <= 0;
        retro_main_state <= retro_main_L3_while432_S3;
      end
      retro_main_L3_while432_S3: begin
        /* cmd_reply_inl2_inl1_inl51 <= (t983_inl2_inl1_inl51 & 4294967295); */
        /* c985_inl2_inl1_inl51 <= (cmd_reply_inl2_inl1_inl51 == 2147483650); */
        if (c985_inl2_inl1_inl51) begin
          io_ports_addr <= 3;
          io_ports_we <= 0;
          io_ports_req <= 1;
          retro_main_state <= retro_main_L1_whileexit434_S1;
        end else begin
          /* c2907 <= (c2901 && !c985_inl2_inl1_inl51); */
          /* c2283 <= (c2243 && !c985_inl2_inl1_inl51); */
          retro_main_state <= retro_main_L3_while432_S0;
        end
      end
      retro_main_L4_while437_S0: begin
        io_ports_addr <= 1;
        io_ports_we <= 0;
        io_ports_req <= 1;
        retro_main_state <= retro_main_L4_while437_S1;
      end
      retro_main_L4_while437_S1: begin
        /*wait for output of io_ports*/
        retro_main_state <= retro_main_L4_while437_S2;
      end
      retro_main_L4_while437_S2: begin
        t983_inl3_inl1_inl51 <= io_ports_q;
        io_ports_req <= 0;
        retro_main_state <= retro_main_L4_while437_S3;
      end
      retro_main_L4_while437_S3: begin
        /* cmd_reply_inl3_inl1_inl51 <= (t983_inl3_inl1_inl51 & 4294967295); */
        /* c985_inl3_inl1_inl51 <= (cmd_reply_inl3_inl1_inl51 == 2147483648); */
        if (c985_inl3_inl1_inl51) begin
          array998[1] <= char_c_inl1_inl51;
          retro_main_state <= retro_main_L1_whileexit439_S1;
        end else begin
          /* c2911 <= (c2901 && !c985_inl3_inl1_inl51); */
          /* c2287 <= (c2243 && !c985_inl3_inl1_inl51); */
          retro_main_state <= retro_main_L4_while437_S0;
        end
      end
      retro_main_L5_while576_S0: begin
        io_ports_addr <= 0;
        io_ports_we <= 0;
        io_ports_req <= 1;
        retro_main_state <= retro_main_L5_while576_S1;
      end
      retro_main_L5_while576_S1: begin
        /*wait for output of io_ports*/
        retro_main_state <= retro_main_L5_while576_S2;
      end
      retro_main_L5_while576_S2: begin
        t992_inl1_inl8_inl51 <= io_ports_q;
        io_ports_req <= 0;
        retro_main_state <= retro_main_L5_while576_S3;
      end
      retro_main_L5_while576_S3: begin
        /* cmd_reply_inl1_inl8_inl51 <= (t992_inl1_inl8_inl51 & 4294967295); */
        /* t993_inl1_inl8_inl51 <= (cmd_reply_inl1_inl8_inl51 & 2147483648); */
        /* c994_inl1_inl8_inl51 <= (t993_inl1_inl8_inl51 == 0); */
        if (c994_inl1_inl8_inl51) begin
          io_ports_addr <= 3;
          io_ports_we <= 1;
          io_ports_req <= 1;
          io_ports_d <= stack0_top2;
          retro_main_state <= retro_main_L1_whileexit578_S1;
        end else begin
          /* c2922 <= (c2920 && !c994_inl1_inl8_inl51); */
          /* c2311 <= (c2301 && !c994_inl1_inl8_inl51); */
          retro_main_state <= retro_main_L5_while576_S0;
        end
      end
      retro_main_L6_while581_S0: begin
        io_ports_addr <= 1;
        io_ports_we <= 0;
        io_ports_req <= 1;
        retro_main_state <= retro_main_L6_while581_S1;
      end
      retro_main_L6_while581_S1: begin
        /*wait for output of io_ports*/
        retro_main_state <= retro_main_L6_while581_S2;
      end
      retro_main_L6_while581_S2: begin
        t983_inl2_inl8_inl51 <= io_ports_q;
        io_ports_req <= 0;
        retro_main_state <= retro_main_L6_while581_S3;
      end
      retro_main_L6_while581_S3: begin
        /* cmd_reply_inl2_inl8_inl51 <= (t983_inl2_inl8_inl51 & 4294967295); */
        /* c985_inl2_inl8_inl51 <= (cmd_reply_inl2_inl8_inl51 == 2147483649); */
        if (c985_inl2_inl8_inl51) begin
          io_ports_addr <= 1;
          io_ports_we <= 1;
          io_ports_req <= 1;
          io_ports_d <= 0;
          retro_main_state <= retro_main_L1_whileexit583_S1;
        end else begin
          /* c2924 <= (c2920 && !c985_inl2_inl8_inl51); */
          /* c2313 <= (c2301 && !c985_inl2_inl8_inl51); */
          retro_main_state <= retro_main_L6_while581_S0;
        end
      end
      retro_main_L7_while586_S0: begin
        io_ports_addr <= 1;
        io_ports_we <= 0;
        io_ports_req <= 1;
        retro_main_state <= retro_main_L7_while586_S1;
      end
      retro_main_L7_while586_S1: begin
        /*wait for output of io_ports*/
        retro_main_state <= retro_main_L7_while586_S2;
      end
      retro_main_L7_while586_S2: begin
        t983_inl3_inl8_inl51 <= io_ports_q;
        io_ports_req <= 0;
        retro_main_state <= retro_main_L7_while586_S3;
      end
      retro_main_L7_while586_S3: begin
        /* cmd_reply_inl3_inl8_inl51 <= (t983_inl3_inl8_inl51 & 4294967295); */
        /* c985_inl3_inl8_inl51 <= (cmd_reply_inl3_inl8_inl51 == 2147483648); */
        if (c985_inl3_inl8_inl51) begin
          /* stack0_pos33 <= (c2300 && c985_inl3_inl7_inl51) ? stack0_pos30 : (c2301 && c985_inl3_inl8_inl51) ? stack0_pos31 : c2298 ? stack0_pos32 : 'bz; */
          /* c2932 <= (c2920 && c985_inl3_inl8_inl51); */
          /* c2933 <= (c2919 && c985_inl3_inl7_inl51); */
          /* stack0_second35 <= (c2300 && c985_inl3_inl7_inl51) ? stack0_second32 : (c2301 && c985_inl3_inl8_inl51) ? stack0_second33 : c2298 ? stack0_second34 : 'bz; */
          /* c2322 <= (c2301 && c985_inl3_inl8_inl51); */
          /* c2323 <= (c2300 && c985_inl3_inl7_inl51); */
          retro_main_state <= retro_main_L17_while505_S0;
        end else begin
          /* c2926 <= (c2920 && !c985_inl3_inl8_inl51); */
          /* c2315 <= (c2301 && !c985_inl3_inl8_inl51); */
          retro_main_state <= retro_main_L7_while586_S0;
        end
      end
      retro_main_L8_while453_S0: begin
        io_ports_addr <= 0;
        io_ports_we <= 0;
        io_ports_req <= 1;
        retro_main_state <= retro_main_L8_while453_S1;
      end
      retro_main_L8_while453_S1: begin
        /*wait for output of io_ports*/
        retro_main_state <= retro_main_L8_while453_S2;
      end
      retro_main_L8_while453_S2: begin
        t992_inl1_inl5_inl51 <= io_ports_q;
        io_ports_req <= 0;
        retro_main_state <= retro_main_L8_while453_S3;
      end
      retro_main_L8_while453_S3: begin
        /* cmd_reply_inl1_inl5_inl51 <= (t992_inl1_inl5_inl51 & 4294967295); */
        /* t993_inl1_inl5_inl51 <= (cmd_reply_inl1_inl5_inl51 & 2147483648); */
        /* c994_inl1_inl5_inl51 <= (t993_inl1_inl5_inl51 == 0); */
        if (c994_inl1_inl5_inl51) begin
          io_ports_addr <= 3;
          io_ports_we <= 1;
          io_ports_req <= 1;
          io_ports_d <= stack0_top2;
          retro_main_state <= retro_main_L1_whileexit455_S1;
        end else begin
          /* c2921 <= (c2919 && !c994_inl1_inl5_inl51); */
          /* c2310 <= (c2300 && !c994_inl1_inl5_inl51); */
          retro_main_state <= retro_main_L8_while453_S0;
        end
      end
      retro_main_L9_while458_S0: begin
        io_ports_addr <= 1;
        io_ports_we <= 0;
        io_ports_req <= 1;
        retro_main_state <= retro_main_L9_while458_S1;
      end
      retro_main_L9_while458_S1: begin
        /*wait for output of io_ports*/
        retro_main_state <= retro_main_L9_while458_S2;
      end
      retro_main_L9_while458_S2: begin
        t983_inl2_inl5_inl51 <= io_ports_q;
        io_ports_req <= 0;
        retro_main_state <= retro_main_L9_while458_S3;
      end
      retro_main_L9_while458_S3: begin
        /* cmd_reply_inl2_inl5_inl51 <= (t983_inl2_inl5_inl51 & 4294967295); */
        /* c985_inl2_inl5_inl51 <= (cmd_reply_inl2_inl5_inl51 == 2147483649); */
        if (c985_inl2_inl5_inl51) begin
          io_ports_addr <= 1;
          io_ports_we <= 1;
          io_ports_req <= 1;
          io_ports_d <= 0;
          retro_main_state <= retro_main_L1_whileexit460_S1;
        end else begin
          /* c2923 <= (c2919 && !c985_inl2_inl5_inl51); */
          /* c2312 <= (c2300 && !c985_inl2_inl5_inl51); */
          retro_main_state <= retro_main_L9_while458_S0;
        end
      end
      endcase
    end
  end
  

endmodule

