module test
  (
    
  );

  //localparams
  localparam CLK_PERIOD = 10;
  localparam CLK_HALF_PERIOD = 5;
  localparam INITIAL_RESET_SPAN = 100;
  localparam test_b1_INIT = 0;
  localparam test_b1_S1 = 1;
  localparam test_b1_S2 = 2;
  localparam test_b1_S3 = 3;
  localparam test_b1_S4 = 4;
  localparam test_b1_S5 = 5;
  localparam test_b1_S6 = 6;
  localparam test_b1_S7 = 7;
  localparam test_b1_S8 = 8;
  localparam test_b1_S9 = 9;
  localparam test_b1_S10 = 10;
  localparam test_b1_S11 = 11;
  localparam test_b1_S12 = 12;
  localparam test_b1_S13 = 13;
  localparam test_b1_S14 = 14;
  localparam test_b1_S15 = 15;
  localparam test_b1_S16 = 16;
  localparam test_b1_S17 = 17;
  localparam test_b1_S18 = 18;
  localparam test_b1_S19 = 19;
  localparam test_b1_S20 = 20;
  localparam test_b1_S21 = 21;
  localparam test_b1_S22 = 22;
  localparam test_b1_S23 = 23;
  localparam test_b1_S24 = 24;
  localparam test_b1_S25 = 25;
  localparam test_b1_S26 = 26;
  localparam test_b1_S27 = 27;
  localparam test_b1_S28 = 28;
  localparam test_b1_S29 = 29;
  localparam test_b1_S30 = 30;
  localparam test_b1_S31 = 31;
  localparam test_b1_S32 = 32;
  localparam test_b1_S33 = 33;
  localparam test_b1_S34 = 34;
  localparam test_b1_S35 = 35;
  localparam test_b1_S36 = 36;
  localparam test_b1_S37 = 37;
  localparam test_b1_S38 = 38;
  localparam test_b1_S39 = 39;
  localparam test_b1_S40 = 40;
  localparam test_b1_S41 = 41;
  localparam test_b1_S42 = 42;
  localparam test_b1_S43 = 43;
  localparam test_b1_S44 = 44;
  localparam test_b1_S45 = 45;
  localparam test_b1_S46 = 46;
  localparam test_b1_S47 = 47;
  localparam test_b1_S48 = 48;
  localparam test_b1_S49 = 49;
  localparam test_b1_S50 = 50;
  localparam test_b1_S51 = 51;
  localparam test_b1_S52 = 52;
  localparam test_b1_S53 = 53;
  localparam test_b1_S54 = 54;
  localparam test_b1_S55 = 55;
  localparam test_b1_S56 = 56;
  localparam test_b1_S57 = 57;
  localparam test_b1_S58 = 58;
  localparam test_b1_S59 = 59;
  localparam test_b1_S60 = 60;
  localparam test_b1_S61 = 61;
  localparam test_b1_S62 = 62;
  localparam test_b1_S63 = 63;
  localparam test_b1_S64 = 64;
  localparam test_b1_S65 = 65;
  localparam test_b1_S66 = 66;
  localparam test_b1_S67 = 67;
  localparam test_b1_S68 = 68;
  localparam test_b1_S69 = 69;
  localparam test_b1_S70 = 70;
  localparam test_b1_S71 = 71;
  localparam test_b1_S72 = 72;
  localparam test_b1_S73 = 73;
  localparam test_b1_S74 = 74;
  localparam test_b1_S75 = 75;
  localparam test_b1_S76 = 76;
  localparam test_b1_S77 = 77;
  localparam test_b1_S78 = 78;
  localparam test_b1_S79 = 79;
  localparam test_b1_S80 = 80;
  localparam test_b1_S81 = 81;
  localparam test_b1_S82 = 82;
  localparam test_b1_S83 = 83;
  localparam test_b1_S84 = 84;
  localparam test_b1_S85 = 85;
  localparam test_b1_S86 = 86;
  localparam test_b1_S87 = 87;
  localparam test_b1_S88 = 88;
  localparam test_b1_S89 = 89;
  localparam test_b1_S90 = 90;
  localparam test_b1_S91 = 91;
  localparam test_b1_S92 = 92;
  localparam test_b1_S93 = 93;
  localparam test_b1_S94 = 94;
  localparam test_b1_S95 = 95;
  localparam test_b1_S96 = 96;
  localparam test_b1_S97 = 97;
  localparam test_b1_S98 = 98;
  localparam test_b1_S99 = 99;
  localparam test_b1_S100 = 100;
  localparam test_b1_S101 = 101;
  localparam test_b1_S102 = 102;
  localparam test_b1_S103 = 103;
  localparam test_b1_S104 = 104;
  localparam test_b1_S105 = 105;
  localparam test_b1_S106 = 106;
  localparam test_b1_S107 = 107;
  localparam test_b1_S108 = 108;
  localparam test_b1_S109 = 109;
  localparam test_b1_S110 = 110;
  localparam test_b1_S111 = 111;
  localparam test_b1_S112 = 112;
  localparam test_b1_S113 = 113;
  localparam test_b1_S114 = 114;
  localparam test_b1_S115 = 115;
  localparam test_b1_S116 = 116;
  localparam test_b1_S117 = 117;
  localparam test_b1_S118 = 118;
  localparam test_b1_S119 = 119;
  localparam test_b1_S120 = 120;
  localparam test_b1_S121 = 121;
  localparam test_b1_S122 = 122;
  localparam test_b1_S123 = 123;
  localparam test_b1_S124 = 124;
  localparam test_b1_S125 = 125;
  localparam test_b1_S126 = 126;
  localparam test_b1_S127 = 127;
  localparam test_b1_S128 = 128;
  localparam test_b1_S129 = 129;
  localparam test_b1_S130 = 130;
  localparam test_b1_S131 = 131;
  localparam test_b1_S132 = 132;
  localparam test_b1_S133 = 133;
  localparam test_b1_S134 = 134;
  localparam test_b1_S135 = 135;
  localparam test_b1_S136 = 136;
  localparam test_b1_S137 = 137;
  localparam test_b1_S138 = 138;
  localparam test_b1_S139 = 139;
  localparam test_b1_S140 = 140;
  localparam test_b1_S141 = 141;
  localparam test_b1_S142 = 142;
  localparam test_b1_S143 = 143;
  localparam test_b1_S144 = 144;
  localparam test_b1_S145 = 145;
  localparam test_b1_S146 = 146;
  localparam test_b1_S147 = 147;
  localparam test_b1_S148 = 148;
  localparam test_b1_S149 = 149;
  localparam test_b1_S150 = 150;
  localparam test_b1_S151 = 151;
  localparam test_b1_S152 = 152;
  localparam test_b1_S153 = 153;
  localparam test_b1_S154 = 154;
  localparam test_b1_S155 = 155;
  localparam test_b1_S156 = 156;
  localparam test_b1_S157 = 157;
  localparam test_b1_S158 = 158;
  localparam test_b1_S159 = 159;
  localparam test_b1_S160 = 160;
  localparam test_b1_S161 = 161;
  localparam test_b1_S162 = 162;
  localparam test_b1_S163 = 163;
  localparam test_b1_S164 = 164;
  localparam test_b1_S165 = 165;
  localparam test_b1_S166 = 166;
  localparam test_b1_S167 = 167;
  localparam test_b1_S168 = 168;
  localparam test_b1_S169 = 169;
  localparam test_b1_S170 = 170;
  localparam test_b1_S171 = 171;
  localparam test_b1_S172 = 172;
  localparam test_b1_S173 = 173;
  localparam test_b1_S174 = 174;
  localparam test_b1_S175 = 175;
  localparam test_b1_S176 = 176;
  localparam test_b1_S177 = 177;
  localparam test_b1_S178 = 178;
  localparam test_b1_S179 = 179;
  localparam test_b1_S180 = 180;
  localparam test_b1_S181 = 181;
  localparam test_b1_S182 = 182;
  localparam test_b1_S183 = 183;
  localparam test_b1_S184 = 184;
  localparam test_b1_S185 = 185;
  localparam test_b1_S186 = 186;
  localparam test_b1_S187 = 187;
  localparam test_b1_S188 = 188;
  localparam test_b1_S189 = 189;
  localparam test_b1_S190 = 190;
  localparam test_b1_S191 = 191;
  localparam test_b1_S192 = 192;
  localparam test_b1_S193 = 193;
  localparam test_b1_S194 = 194;
  localparam test_b1_S195 = 195;
  localparam test_b1_S196 = 196;
  localparam test_b1_S197 = 197;
  localparam test_b1_S198 = 198;
  localparam test_b1_S199 = 199;
  localparam test_b1_S200 = 200;
  localparam test_b1_S201 = 201;
  localparam test_b1_S202 = 202;
  localparam test_b1_S203 = 203;
  localparam test_b1_S204 = 204;
  localparam test_b1_S205 = 205;
  localparam test_b1_S206 = 206;
  localparam test_b1_S207 = 207;
  localparam test_b1_S208 = 208;
  localparam test_b1_S209 = 209;
  localparam test_b1_S210 = 210;
  localparam test_b1_S211 = 211;
  localparam test_b1_S212 = 212;
  localparam test_b1_S213 = 213;
  localparam test_b1_S214 = 214;
  localparam test_b1_S215 = 215;
  localparam test_b1_S216 = 216;
  localparam test_b1_S217 = 217;
  localparam test_b1_S218 = 218;
  localparam test_b1_S219 = 219;
  localparam test_b1_S220 = 220;
  localparam test_b1_S221 = 221;
  localparam test_b1_S222 = 222;
  localparam test_b1_S223 = 223;
  localparam test_b1_S224 = 224;
  localparam test_b1_S225 = 225;
  localparam test_b1_S226 = 226;
  localparam test_b1_S227 = 227;
  localparam test_b1_S228 = 228;
  localparam test_b1_S229 = 229;
  localparam test_b1_S230 = 230;
  localparam test_b1_S231 = 231;
  localparam test_b1_S232 = 232;
  localparam test_b1_S233 = 233;
  localparam test_b1_S234 = 234;
  localparam test_b1_S235 = 235;
  localparam test_b1_S236 = 236;
  localparam test_b1_S237 = 237;
  localparam test_b1_S238 = 238;
  localparam test_b1_S239 = 239;
  localparam test_b1_S240 = 240;
  localparam test_b1_S241 = 241;
  localparam test_b1_S242 = 242;
  localparam test_b1_S243 = 243;
  localparam test_b1_S244 = 244;
  localparam test_b1_S245 = 245;
  localparam test_b1_S246 = 246;
  localparam test_b1_S247 = 247;
  localparam test_b1_S248 = 248;
  localparam test_b1_S249 = 249;
  localparam test_b1_S250 = 250;
  localparam test_b1_S251 = 251;
  localparam test_b1_S252 = 252;
  localparam test_b1_S253 = 253;
  localparam test_b1_S254 = 254;
  localparam test_b1_S255 = 255;
  localparam test_b1_S256 = 256;
  localparam test_b1_S257 = 257;
  localparam test_b1_S258 = 258;
  localparam test_b1_S259 = 259;
  localparam test_b1_S260 = 260;
  localparam test_b1_S261 = 261;
  localparam test_b1_S262 = 262;
  localparam test_b1_S263 = 263;
  localparam test_b1_S264 = 264;
  localparam test_b1_S265 = 265;
  localparam test_b1_S266 = 266;
  localparam test_b1_S267 = 267;
  localparam test_b1_S268 = 268;
  localparam test_b1_S269 = 269;
  localparam test_b1_S270 = 270;
  localparam test_b1_S271 = 271;
  localparam test_b1_S272 = 272;
  localparam test_b1_S273 = 273;
  localparam test_b1_S274 = 274;
  localparam test_b1_S275 = 275;
  localparam test_b1_S276 = 276;
  localparam test_b1_S277 = 277;
  localparam test_b1_S278 = 278;
  localparam test_b1_S279 = 279;
  localparam test_b1_S280 = 280;
  localparam test_b1_S281 = 281;
  localparam test_b1_S282 = 282;
  localparam test_b1_S283 = 283;
  localparam test_b1_S284 = 284;
  localparam test_b1_S285 = 285;
  localparam test_b1_S286 = 286;
  localparam test_b1_S287 = 287;
  localparam test_b1_S288 = 288;
  localparam test_b1_S289 = 289;
  localparam test_b1_S290 = 290;
  localparam test_b1_S291 = 291;
  localparam test_b1_S292 = 292;
  localparam test_b1_S293 = 293;
  localparam test_b1_S294 = 294;
  localparam test_b1_S295 = 295;
  localparam test_b1_S296 = 296;
  localparam test_b1_S297 = 297;
  localparam test_b1_S298 = 298;
  localparam test_b1_S299 = 299;
  localparam test_b1_S300 = 300;
  localparam test_b1_S301 = 301;
  localparam test_b1_S302 = 302;
  localparam test_b1_S303 = 303;
  localparam test_b1_S304 = 304;
  localparam test_b1_S305 = 305;
  localparam test_b1_S306 = 306;
  localparam test_b1_S307 = 307;
  localparam test_b1_S308 = 308;
  localparam test_b1_S309 = 309;
  localparam test_b1_S310 = 310;
  localparam test_b1_S311 = 311;
  localparam test_b1_S312 = 312;
  localparam test_b1_S313 = 313;
  localparam test_b1_S314 = 314;
  localparam test_b1_S315 = 315;
  localparam test_b1_S316 = 316;
  localparam test_b1_S317 = 317;
  localparam test_b1_S318 = 318;
  localparam test_b1_S319 = 319;
  localparam test_b1_S320 = 320;
  localparam test_b1_S321 = 321;
  localparam test_b1_S322 = 322;
  localparam test_b1_S323 = 323;
  localparam test_b1_S324 = 324;
  localparam test_b1_S325 = 325;
  localparam test_b1_S326 = 326;
  localparam test_b1_S327 = 327;
  localparam test_b1_S328 = 328;
  localparam test_b1_S329 = 329;
  localparam test_b1_S330 = 330;
  localparam test_b1_S331 = 331;
  localparam test_b1_S332 = 332;
  localparam test_b1_S333 = 333;
  localparam test_b1_S334 = 334;
  localparam test_b1_S335 = 335;
  localparam test_b1_S336 = 336;
  localparam test_b1_S337 = 337;
  localparam test_b1_S338 = 338;
  localparam test_b1_S339 = 339;
  localparam test_b1_S340 = 340;
  localparam test_b1_S341 = 341;
  localparam test_b1_S342 = 342;
  localparam test_b1_S343 = 343;
  localparam test_b1_S344 = 344;
  localparam test_b1_S345 = 345;
  localparam test_b1_S346 = 346;
  localparam test_b1_S347 = 347;
  localparam test_b1_S348 = 348;
  localparam test_b1_S349 = 349;
  localparam test_b1_S350 = 350;
  localparam test_b1_S351 = 351;
  localparam test_b1_S352 = 352;
  localparam test_b1_S353 = 353;
  localparam test_b1_S354 = 354;
  localparam test_b1_S355 = 355;
  localparam test_b1_S356 = 356;
  localparam test_b1_S357 = 357;
  localparam test_b1_S358 = 358;
  localparam test_b1_S359 = 359;
  localparam test_b1_S360 = 360;
  localparam test_b1_S361 = 361;
  localparam test_b1_S362 = 362;
  localparam test_b1_S363 = 363;
  localparam test_b1_S364 = 364;
  localparam test_b1_S365 = 365;
  localparam test_b1_S366 = 366;
  localparam test_b1_S367 = 367;
  localparam test_b1_S368 = 368;
  localparam test_b1_S369 = 369;
  localparam test_b1_S370 = 370;
  localparam test_b1_S371 = 371;
  localparam test_b1_S372 = 372;
  localparam test_b1_S373 = 373;
  localparam test_b1_S374 = 374;
  localparam test_b1_S375 = 375;
  localparam test_b1_S376 = 376;
  localparam test_b1_S377 = 377;
  localparam test_b1_S378 = 378;
  localparam test_b1_S379 = 379;
  localparam test_b1_S380 = 380;
  localparam test_b1_S381 = 381;
  localparam test_b1_S382 = 382;
  localparam test_b1_S383 = 383;
  localparam test_b1_S384 = 384;
  localparam test_b1_S385 = 385;
  localparam test_b1_S386 = 386;
  localparam test_b1_S387 = 387;
  localparam test_b1_S388 = 388;
  localparam test_b1_S389 = 389;
  localparam test_b1_S390 = 390;
  localparam test_b1_S391 = 391;
  localparam test_b1_S392 = 392;
  localparam test_b1_S393 = 393;
  localparam test_b1_S394 = 394;
  localparam test_b1_S395 = 395;
  localparam test_b1_S396 = 396;
  localparam test_b1_S397 = 397;
  localparam test_b1_S398 = 398;
  localparam test_b1_S399 = 399;
  localparam test_b1_S400 = 400;
  localparam test_b1_S401 = 401;
  localparam test_b1_S402 = 402;
  localparam test_b1_S403 = 403;
  localparam test_b1_S404 = 404;
  localparam test_b1_S405 = 405;
  localparam test_b1_S406 = 406;
  localparam test_b1_S407 = 407;
  localparam test_b1_S408 = 408;
  localparam test_b1_S409 = 409;
  localparam test_b1_S410 = 410;
  localparam test_b1_S411 = 411;
  localparam test_b1_S412 = 412;
  localparam test_b1_S413 = 413;
  localparam test_b1_S414 = 414;
  localparam test_b1_S415 = 415;
  localparam test_b1_S416 = 416;
  localparam test_b1_S417 = 417;
  localparam test_b1_S418 = 418;
  localparam test_b1_S419 = 419;
  localparam test_b1_S420 = 420;
  localparam test_b1_S421 = 421;
  localparam test_b1_S422 = 422;
  localparam test_b1_S423 = 423;
  localparam test_b1_S424 = 424;
  localparam test_b1_S425 = 425;
  localparam test_b1_S426 = 426;
  localparam test_b1_S427 = 427;
  localparam test_b1_S428 = 428;
  localparam test_b1_S429 = 429;
  localparam test_b1_S430 = 430;
  localparam test_b1_S431 = 431;
  localparam test_b1_S432 = 432;
  localparam test_b1_S433 = 433;
  localparam test_b1_S434 = 434;
  localparam test_b1_S435 = 435;
  localparam test_b1_S436 = 436;
  localparam test_b1_S437 = 437;
  localparam test_b1_S438 = 438;
  localparam test_b1_S439 = 439;
  localparam test_b1_S440 = 440;
  localparam test_b1_S441 = 441;
  localparam test_b1_S442 = 442;
  localparam test_b1_S443 = 443;
  localparam test_b1_S444 = 444;
  localparam test_b1_S445 = 445;
  localparam test_b1_S446 = 446;
  localparam test_b1_S447 = 447;
  localparam test_b1_S448 = 448;
  localparam test_b1_S449 = 449;
  localparam test_b1_S450 = 450;
  localparam test_b1_S451 = 451;
  localparam test_b1_S452 = 452;
  localparam test_b1_S453 = 453;
  localparam test_b1_S454 = 454;
  localparam test_b1_S455 = 455;
  localparam test_b1_S456 = 456;
  localparam test_b1_S457 = 457;
  localparam test_b1_S458 = 458;
  localparam test_b1_S459 = 459;
  localparam test_b1_S460 = 460;
  localparam test_b1_S461 = 461;
  localparam test_b1_S462 = 462;
  localparam test_b1_S463 = 463;
  localparam test_b1_S464 = 464;
  localparam test_b1_S465 = 465;
  localparam test_b1_S466 = 466;
  localparam test_b1_S467 = 467;
  localparam test_b1_S468 = 468;
  localparam test_b1_S469 = 469;
  localparam test_b1_S470 = 470;
  localparam test_b1_S471 = 471;
  localparam test_b1_S472 = 472;
  localparam test_b1_S473 = 473;
  localparam test_b1_S474 = 474;
  localparam test_b1_S475 = 475;
  localparam test_b1_S476 = 476;
  localparam test_b1_S477 = 477;
  localparam test_b1_S478 = 478;
  localparam test_b1_S479 = 479;
  localparam test_b1_S480 = 480;
  localparam test_b1_S481 = 481;
  localparam test_b1_S482 = 482;
  localparam test_b1_S483 = 483;
  localparam test_b1_S484 = 484;
  localparam test_b1_S485 = 485;
  localparam test_b1_S486 = 486;
  localparam test_b1_S487 = 487;
  localparam test_b1_S488 = 488;
  localparam test_b1_S489 = 489;
  localparam test_b1_S490 = 490;
  localparam test_b1_S491 = 491;
  localparam test_b1_S492 = 492;
  localparam test_b1_S493 = 493;
  localparam test_b1_S494 = 494;
  localparam test_b1_S495 = 495;
  localparam test_b1_S496 = 496;
  localparam test_b1_S497 = 497;
  localparam test_b1_S498 = 498;
  localparam test_b1_S499 = 499;
  localparam test_b1_S500 = 500;
  localparam test_b1_S501 = 501;
  localparam test_b1_S502 = 502;
  localparam test_b1_S503 = 503;
  localparam test_b1_S504 = 504;
  localparam test_b1_S505 = 505;
  localparam test_b1_S506 = 506;
  localparam test_b1_S507 = 507;
  localparam test_b1_S508 = 508;
  localparam test_b1_S509 = 509;
  localparam test_b1_S510 = 510;
  localparam test_b1_S511 = 511;
  localparam test_b1_S512 = 512;
  localparam test_b1_S513 = 513;
  localparam test_b1_S514 = 514;
  localparam test_b1_S515 = 515;
  localparam test_b1_S516 = 516;
  localparam test_b1_S517 = 517;
  localparam test_b1_S518 = 518;
  localparam test_b1_S519 = 519;
  localparam test_b1_S520 = 520;
  localparam test_b1_S521 = 521;
  localparam test_b1_S522 = 522;
  localparam test_b1_S523 = 523;
  localparam test_b1_S524 = 524;
  localparam test_b1_S525 = 525;
  localparam test_b1_S526 = 526;
  localparam test_b1_S527 = 527;
  localparam test_b1_S528 = 528;
  localparam test_b1_S529 = 529;
  localparam test_b1_S530 = 530;
  localparam test_b1_S531 = 531;
  localparam test_b1_S532 = 532;
  localparam test_b1_S533 = 533;
  localparam test_b1_S534 = 534;
  localparam test_b1_S535 = 535;
  localparam test_b1_S536 = 536;
  localparam test_b1_S537 = 537;
  localparam test_b1_S538 = 538;
  localparam test_b1_S539 = 539;
  localparam test_b1_S540 = 540;
  localparam test_b1_S541 = 541;
  localparam test_b1_S542 = 542;
  localparam test_b1_S543 = 543;
  localparam test_b1_S544 = 544;
  localparam test_b1_S545 = 545;
  localparam test_b1_S546 = 546;
  localparam test_b1_S547 = 547;
  localparam test_b1_S548 = 548;
  localparam test_b1_S549 = 549;
  localparam test_b1_S550 = 550;
  localparam test_b1_S551 = 551;
  localparam test_b1_S552 = 552;
  localparam test_b1_S553 = 553;
  localparam test_b1_S554 = 554;
  localparam test_b1_S555 = 555;
  localparam test_b1_S556 = 556;
  localparam test_b1_S557 = 557;
  localparam test_b1_S558 = 558;
  localparam test_b1_S559 = 559;
  localparam test_b1_S560 = 560;
  localparam test_b1_S561 = 561;
  localparam test_b1_S562 = 562;
  localparam test_b1_S563 = 563;
  localparam test_b1_S564 = 564;
  localparam test_b1_S565 = 565;
  localparam test_b1_S566 = 566;
  localparam test_b1_S567 = 567;
  localparam test_b1_S568 = 568;
  localparam test_b1_S569 = 569;
  localparam test_b1_S570 = 570;
  localparam test_b1_S571 = 571;
  localparam test_b1_S572 = 572;
  localparam test_b1_S573 = 573;
  localparam test_b1_S574 = 574;
  localparam test_b1_S575 = 575;
  localparam test_b1_S576 = 576;
  localparam test_b1_S577 = 577;
  localparam test_b1_S578 = 578;
  localparam test_b1_S579 = 579;
  localparam test_b1_S580 = 580;
  localparam test_b1_S581 = 581;
  localparam test_b1_S582 = 582;
  localparam test_b1_S583 = 583;
  localparam test_b1_S584 = 584;
  localparam test_b1_S585 = 585;
  localparam test_b1_S586 = 586;
  localparam test_b1_S587 = 587;
  localparam test_b1_S588 = 588;
  localparam test_b1_S589 = 589;
  localparam test_b1_S590 = 590;
  localparam test_b1_S591 = 591;
  localparam test_b1_S592 = 592;
  localparam test_b1_S593 = 593;
  localparam test_b1_S594 = 594;
  localparam test_b1_S595 = 595;
  localparam test_b1_S596 = 596;
  localparam test_b1_S597 = 597;
  localparam test_b1_S598 = 598;
  localparam test_b1_S599 = 599;
  localparam test_b1_S600 = 600;
  localparam test_b1_S601 = 601;
  localparam test_b1_S602 = 602;
  localparam test_b1_S603 = 603;
  localparam test_b1_S604 = 604;
  localparam test_b1_S605 = 605;
  localparam test_b1_S606 = 606;
  localparam test_b1_S607 = 607;
  localparam test_b1_S608 = 608;
  localparam test_b1_S609 = 609;
  localparam test_b1_S610 = 610;
  localparam test_b1_S611 = 611;
  localparam test_b1_S612 = 612;
  localparam test_b1_S613 = 613;
  localparam test_b1_S614 = 614;
  localparam test_b1_S615 = 615;
  localparam test_b1_S616 = 616;
  localparam test_b1_S617 = 617;
  localparam test_b1_S618 = 618;
  localparam test_b1_S619 = 619;
  localparam test_b1_S620 = 620;
  localparam test_b1_S621 = 621;
  localparam test_b1_S622 = 622;
  localparam test_b1_S623 = 623;
  localparam test_b1_S624 = 624;
  localparam test_b1_S625 = 625;
  localparam test_b1_S626 = 626;
  localparam test_b1_S627 = 627;
  localparam test_b1_S628 = 628;
  localparam test_b1_S629 = 629;
  localparam test_b1_S630 = 630;
  localparam test_b1_S631 = 631;
  localparam test_b1_S632 = 632;
  localparam test_b1_S633 = 633;
  localparam test_b1_S634 = 634;
  localparam test_b1_S635 = 635;
  localparam test_b1_S636 = 636;
  localparam test_b1_S637 = 637;
  localparam test_b1_S638 = 638;
  localparam test_b1_S639 = 639;
  localparam test_b1_S640 = 640;
  localparam test_b1_S641 = 641;
  localparam test_b1_S642 = 642;
  localparam test_b1_S643 = 643;
  localparam test_b1_S644 = 644;
  localparam test_b1_S645 = 645;
  localparam test_b1_S646 = 646;
  localparam test_b1_S647 = 647;
  localparam test_b1_S648 = 648;
  localparam test_b1_S649 = 649;
  localparam test_b1_S650 = 650;
  localparam test_b1_S651 = 651;
  localparam test_b1_S652 = 652;
  localparam test_b1_S653 = 653;
  localparam test_b1_S654 = 654;
  localparam test_b1_S655 = 655;
  localparam test_b1_S656 = 656;
  localparam test_b1_S657 = 657;
  localparam test_b1_S658 = 658;
  localparam test_b1_S659 = 659;
  localparam test_b1_S660 = 660;
  localparam test_b1_S661 = 661;
  localparam test_b1_S662 = 662;
  localparam test_b1_S663 = 663;
  localparam test_b1_S664 = 664;
  localparam test_b1_S665 = 665;
  localparam test_b1_S666 = 666;
  localparam test_b1_S667 = 667;
  localparam test_b1_S668 = 668;
  localparam test_b1_S669 = 669;
  localparam test_b1_S670 = 670;
  localparam test_b1_S671 = 671;
  localparam test_b1_S672 = 672;
  localparam test_b1_S673 = 673;
  localparam test_b1_S674 = 674;
  localparam test_b1_S675 = 675;
  localparam test_b1_S676 = 676;
  localparam test_b1_S677 = 677;
  localparam test_b1_S678 = 678;
  localparam test_b1_S679 = 679;
  localparam test_b1_S680 = 680;
  localparam test_b1_S681 = 681;
  localparam test_b1_S682 = 682;
  localparam test_b1_S683 = 683;
  localparam test_b1_S684 = 684;
  localparam test_b1_S685 = 685;
  localparam test_b1_S686 = 686;
  localparam test_b1_S687 = 687;
  localparam test_b1_S688 = 688;
  localparam test_b1_S689 = 689;
  localparam test_b1_S690 = 690;
  localparam test_b1_S691 = 691;
  localparam test_b1_S692 = 692;
  localparam test_b1_S693 = 693;
  localparam test_b1_S694 = 694;
  localparam test_b1_S695 = 695;
  localparam test_b1_S696 = 696;
  localparam test_b1_S697 = 697;
  localparam test_b1_S698 = 698;
  localparam test_b1_S699 = 699;
  localparam test_b1_S700 = 700;
  localparam test_b1_S701 = 701;
  localparam test_b1_S702 = 702;
  localparam test_b1_S703 = 703;
  localparam test_b1_S704 = 704;
  localparam test_b1_S705 = 705;
  localparam test_b1_S706 = 706;
  localparam test_b1_S707 = 707;
  localparam test_b1_S708 = 708;
  localparam test_b1_S709 = 709;
  localparam test_b1_S710 = 710;
  localparam test_b1_S711 = 711;
  localparam test_b1_S712 = 712;
  localparam test_b1_S713 = 713;
  localparam test_b1_S714 = 714;
  localparam test_b1_S715 = 715;
  localparam test_b1_S716 = 716;
  localparam test_b1_S717 = 717;
  localparam test_b1_S718 = 718;
  localparam test_b1_S719 = 719;
  localparam test_b1_S720 = 720;
  localparam test_b1_S721 = 721;
  localparam test_b1_S722 = 722;
  localparam test_b1_S723 = 723;
  localparam test_b1_S724 = 724;
  localparam test_b1_S725 = 725;
  localparam test_b1_S726 = 726;
  localparam test_b1_S727 = 727;
  localparam test_b1_S728 = 728;
  localparam test_b1_S729 = 729;
  localparam test_b1_S730 = 730;
  localparam test_b1_S731 = 731;
  localparam test_b1_S732 = 732;
  localparam test_b1_S733 = 733;
  localparam test_b1_S734 = 734;
  localparam test_b1_S735 = 735;
  localparam test_b1_S736 = 736;
  localparam test_b1_S737 = 737;
  localparam test_b1_S738 = 738;
  localparam test_b1_S739 = 739;
  localparam test_b1_S740 = 740;
  localparam test_b1_S741 = 741;
  localparam test_b1_S742 = 742;
  localparam test_b1_S743 = 743;
  localparam test_b1_S744 = 744;
  localparam test_b1_S745 = 745;
  localparam test_b1_S746 = 746;
  localparam test_b1_S747 = 747;
  localparam test_b1_S748 = 748;
  localparam test_b1_S749 = 749;
  localparam test_b1_S750 = 750;
  localparam test_b1_S751 = 751;
  localparam test_b1_S752 = 752;
  localparam test_b1_S753 = 753;
  localparam test_b1_S754 = 754;
  localparam test_b1_S755 = 755;
  localparam test_b1_S756 = 756;
  localparam test_b1_S757 = 757;
  localparam test_b1_S758 = 758;
  localparam test_b1_S759 = 759;
  localparam test_b1_S760 = 760;
  localparam test_b1_S761 = 761;
  localparam test_b1_S762 = 762;
  localparam test_b1_S763 = 763;
  localparam test_b1_S764 = 764;
  localparam test_b1_S765 = 765;
  localparam test_b1_S766 = 766;
  localparam test_b1_S767 = 767;
  localparam test_b1_S768 = 768;
  localparam test_b1_S769 = 769;
  localparam test_b1_S770 = 770;
  localparam test_b1_S771 = 771;
  localparam test_b1_S772 = 772;
  localparam test_b1_S773 = 773;
  localparam test_b1_S774 = 774;
  localparam test_b1_S775 = 775;
  localparam test_b1_S776 = 776;
  localparam test_b1_S777 = 777;
  localparam test_b1_S778 = 778;
  localparam test_b1_S779 = 779;
  localparam test_b1_S780 = 780;
  localparam test_b1_S781 = 781;
  localparam test_b1_S782 = 782;
  localparam test_b1_S783 = 783;
  localparam test_b1_S784 = 784;
  localparam test_b1_S785 = 785;
  localparam test_b1_S786 = 786;
  localparam test_b1_S787 = 787;
  localparam test_b1_S788 = 788;
  localparam test_b1_S789 = 789;
  localparam test_b1_S790 = 790;
  localparam test_b1_S791 = 791;
  localparam test_b1_S792 = 792;
  localparam test_b1_S793 = 793;
  localparam test_b1_S794 = 794;
  localparam test_b1_S795 = 795;
  localparam test_b1_S796 = 796;
  localparam test_b1_S797 = 797;
  localparam test_b1_S798 = 798;
  localparam test_b1_S799 = 799;
  localparam test_b1_S800 = 800;
  localparam test_b1_S801 = 801;
  localparam test_b1_S802 = 802;
  localparam test_b1_S803 = 803;
  localparam test_b1_S804 = 804;
  localparam test_b1_S805 = 805;
  localparam test_b1_S806 = 806;
  localparam test_b1_S807 = 807;
  localparam test_b1_S808 = 808;
  localparam test_b1_S809 = 809;
  localparam test_b1_S810 = 810;
  localparam test_b1_S811 = 811;
  localparam test_b1_S812 = 812;
  localparam test_b1_S813 = 813;
  localparam test_b1_S814 = 814;
  localparam test_b1_S815 = 815;
  localparam test_b1_S816 = 816;
  localparam test_b1_S817 = 817;
  localparam test_b1_S818 = 818;
  localparam test_b1_S819 = 819;
  localparam test_b1_S820 = 820;
  localparam test_b1_S821 = 821;
  localparam test_b1_S822 = 822;
  localparam test_b1_S823 = 823;
  localparam test_b1_S824 = 824;
  localparam test_b1_S825 = 825;
  localparam test_b1_S826 = 826;
  localparam test_b1_S827 = 827;
  localparam test_b1_S828 = 828;
  localparam test_b1_S829 = 829;
  localparam test_b1_S830 = 830;
  localparam test_b1_S831 = 831;
  localparam test_b1_S832 = 832;
  localparam test_b1_S833 = 833;
  localparam test_b1_S834 = 834;
  localparam test_b1_S835 = 835;
  localparam test_b1_S836 = 836;
  localparam test_b1_S837 = 837;
  localparam test_b1_S838 = 838;
  localparam test_b1_S839 = 839;
  localparam test_b1_S840 = 840;
  localparam test_b1_S841 = 841;
  localparam test_b1_S842 = 842;
  localparam test_b1_S843 = 843;
  localparam test_b1_S844 = 844;
  localparam test_b1_S845 = 845;
  localparam test_b1_S846 = 846;
  localparam test_b1_S847 = 847;
  localparam test_b1_S848 = 848;
  localparam test_b1_S849 = 849;
  localparam test_b1_S850 = 850;
  localparam test_b1_S851 = 851;
  localparam test_b1_S852 = 852;
  localparam test_b1_S853 = 853;
  localparam test_b1_S854 = 854;
  localparam test_b1_S855 = 855;
  localparam test_b1_S856 = 856;
  localparam test_b1_S857 = 857;
  localparam test_b1_S858 = 858;
  localparam test_b1_S859 = 859;
  localparam test_b1_S860 = 860;
  localparam test_b1_S861 = 861;
  localparam test_b1_S862 = 862;
  localparam test_b1_S863 = 863;
  localparam test_b1_S864 = 864;
  localparam test_b1_S865 = 865;
  localparam test_b1_S866 = 866;
  localparam test_b1_S867 = 867;
  localparam test_b1_S868 = 868;
  localparam test_b1_S869 = 869;
  localparam test_b1_S870 = 870;
  localparam test_b1_S871 = 871;
  localparam test_b1_S872 = 872;
  localparam test_b1_S873 = 873;
  localparam test_b1_S874 = 874;
  localparam test_b1_S875 = 875;
  localparam test_b1_S876 = 876;
  localparam test_b1_S877 = 877;
  localparam test_b1_S878 = 878;
  localparam test_b1_S879 = 879;
  localparam test_b1_S880 = 880;
  localparam test_b1_S881 = 881;
  localparam test_b1_S882 = 882;
  localparam test_b1_S883 = 883;
  localparam test_b1_S884 = 884;
  localparam test_b1_S885 = 885;
  localparam test_b1_S886 = 886;
  localparam test_b1_S887 = 887;
  localparam test_b1_S888 = 888;
  localparam test_b1_S889 = 889;
  localparam test_b1_S890 = 890;
  localparam test_b1_S891 = 891;
  localparam test_b1_S892 = 892;
  localparam test_b1_S893 = 893;
  localparam test_b1_S894 = 894;
  localparam test_b1_S895 = 895;
  localparam test_b1_S896 = 896;
  localparam test_b1_S897 = 897;
  localparam test_b1_S898 = 898;
  localparam test_b1_S899 = 899;
  localparam test_b1_S900 = 900;
  localparam test_b1_S901 = 901;
  localparam test_b1_S902 = 902;
  localparam test_b1_S903 = 903;
  localparam test_b1_S904 = 904;
  localparam test_b1_S905 = 905;
  localparam test_b1_S906 = 906;
  localparam test_b1_S907 = 907;
  localparam test_b1_S908 = 908;
  localparam test_b1_S909 = 909;
  localparam test_b1_S910 = 910;
  localparam test_b1_S911 = 911;
  localparam test_b1_S912 = 912;
  localparam test_b1_S913 = 913;
  localparam test_b1_S914 = 914;
  localparam test_b1_S915 = 915;
  localparam test_b1_S916 = 916;
  localparam test_b1_S917 = 917;
  localparam test_b1_S918 = 918;
  localparam test_b1_S919 = 919;
  localparam test_b1_S920 = 920;
  localparam test_b1_S921 = 921;
  localparam test_b1_S922 = 922;
  localparam test_b1_S923 = 923;
  localparam test_b1_S924 = 924;
  localparam test_b1_S925 = 925;
  localparam test_b1_S926 = 926;
  localparam test_b1_S927 = 927;
  localparam test_b1_S928 = 928;
  localparam test_b1_S929 = 929;
  localparam test_b1_S930 = 930;
  localparam test_b1_S931 = 931;
  localparam test_b1_S932 = 932;
  localparam test_b1_S933 = 933;
  localparam test_b1_S934 = 934;
  localparam test_b1_S935 = 935;
  localparam test_b1_S936 = 936;
  localparam test_b1_S937 = 937;
  localparam test_b1_S938 = 938;
  localparam test_b1_S939 = 939;
  localparam test_b1_S940 = 940;
  localparam test_b1_S941 = 941;
  localparam test_b1_S942 = 942;
  localparam test_b1_S943 = 943;
  localparam test_b1_S944 = 944;
  localparam test_b1_S945 = 945;
  localparam test_b1_S946 = 946;
  localparam test_b1_S947 = 947;
  localparam test_b1_S948 = 948;
  localparam test_b1_S949 = 949;
  localparam test_b1_S950 = 950;
  localparam test_b1_S951 = 951;
  localparam test_b1_S952 = 952;
  localparam test_b1_S953 = 953;
  localparam test_b1_S954 = 954;
  localparam test_b1_S955 = 955;
  localparam test_b1_S956 = 956;
  localparam test_b1_S957 = 957;
  localparam test_b1_S958 = 958;
  localparam test_b1_S959 = 959;
  localparam test_b1_S960 = 960;
  localparam test_b1_S961 = 961;
  localparam test_b1_S962 = 962;
  localparam test_b1_S963 = 963;
  localparam test_b1_S964 = 964;
  localparam test_b1_S965 = 965;
  localparam test_b1_S966 = 966;
  localparam test_b1_S967 = 967;
  localparam test_b1_S968 = 968;
  localparam test_b1_S969 = 969;
  localparam test_b1_S970 = 970;
  localparam test_b1_S971 = 971;
  localparam test_b1_S972 = 972;
  localparam test_b1_S973 = 973;
  localparam test_b1_S974 = 974;
  localparam test_b1_S975 = 975;
  localparam test_b1_S976 = 976;
  localparam test_b1_S977 = 977;
  localparam test_b1_S978 = 978;
  localparam test_b1_S979 = 979;
  localparam test_b1_S980 = 980;
  localparam test_b1_S981 = 981;
  localparam test_b1_S982 = 982;
  localparam test_b1_S983 = 983;
  localparam test_b1_S984 = 984;
  localparam test_b1_S985 = 985;
  localparam test_b1_S986 = 986;
  localparam test_b1_S987 = 987;
  localparam test_b1_S988 = 988;
  localparam test_b1_S989 = 989;
  localparam test_b1_S990 = 990;
  localparam test_b1_S991 = 991;
  localparam test_b1_S992 = 992;
  localparam test_b1_S993 = 993;
  localparam test_b1_S994 = 994;
  localparam test_b1_S995 = 995;
  localparam test_b1_S996 = 996;
  localparam test_b1_S997 = 997;
  localparam test_b1_S998 = 998;
  localparam test_b1_S999 = 999;
  localparam test_b1_S1000 = 1000;
  localparam test_b1_S1001 = 1001;
  localparam test_b1_S1002 = 1002;
  localparam test_b1_S1003 = 1003;
  localparam test_b1_S1004 = 1004;
  localparam test_b1_S1005 = 1005;
  localparam test_b1_S1006 = 1006;
  localparam test_b1_S1007 = 1007;
  localparam test_b1_S1008 = 1008;
  localparam test_b1_S1009 = 1009;
  localparam test_b1_S1010 = 1010;
  localparam test_b1_S1011 = 1011;
  localparam test_b1_S1012 = 1012;
  localparam test_b1_S1013 = 1013;
  localparam test_b1_S1014 = 1014;
  localparam test_b1_S1015 = 1015;
  localparam test_b1_S1016 = 1016;
  localparam test_b1_S1017 = 1017;
  localparam test_b1_S1018 = 1018;
  localparam test_b1_S1019 = 1019;
  localparam test_b1_S1020 = 1020;
  localparam test_b1_S1021 = 1021;
  localparam test_b1_S1022 = 1022;
  localparam test_b1_S1023 = 1023;
  localparam test_b1_S1024 = 1024;
  localparam test_b1_S1025 = 1025;
  localparam test_b1_S1026 = 1026;
  localparam test_b1_S1027 = 1027;
  localparam test_b1_S1028 = 1028;
  localparam test_b1_S1029 = 1029;
  localparam test_b1_S1030 = 1030;
  localparam test_b1_S1031 = 1031;
  localparam test_b1_S1032 = 1032;
  localparam test_b1_S1033 = 1033;
  localparam test_b1_S1034 = 1034;
  localparam test_b1_S1035 = 1035;
  localparam test_b1_S1036 = 1036;
  localparam test_b1_S1037 = 1037;
  localparam test_b1_S1038 = 1038;
  localparam test_b1_S1039 = 1039;
  localparam test_b1_S1040 = 1040;
  localparam test_b1_S1041 = 1041;
  localparam test_b1_S1042 = 1042;
  localparam test_b1_S1043 = 1043;
  localparam test_b1_S1044 = 1044;
  localparam test_b1_S1045 = 1045;
  localparam test_b1_S1046 = 1046;
  localparam test_b1_S1047 = 1047;
  localparam test_b1_S1048 = 1048;
  localparam test_b1_S1049 = 1049;
  localparam test_b1_S1050 = 1050;
  localparam test_b1_S1051 = 1051;
  localparam test_b1_S1052 = 1052;
  localparam test_b1_S1053 = 1053;
  localparam test_b1_S1054 = 1054;
  localparam test_b1_S1055 = 1055;
  localparam test_b1_S1056 = 1056;
  localparam test_b1_S1057 = 1057;
  localparam test_b1_S1058 = 1058;
  localparam test_b1_S1059 = 1059;
  localparam test_b1_S1060 = 1060;
  localparam test_b1_S1061 = 1061;
  localparam test_b1_S1062 = 1062;
  localparam test_b1_S1063 = 1063;
  localparam test_b1_S1064 = 1064;
  localparam test_b1_S1065 = 1065;
  localparam test_b1_S1066 = 1066;
  localparam test_b1_S1067 = 1067;
  localparam test_b1_S1068 = 1068;
  localparam test_b1_S1069 = 1069;
  localparam test_b1_S1070 = 1070;
  localparam test_b1_S1071 = 1071;
  localparam test_b1_S1072 = 1072;
  localparam test_b1_S1073 = 1073;
  localparam test_b1_S1074 = 1074;
  localparam test_b1_S1075 = 1075;
  localparam test_b1_S1076 = 1076;
  localparam test_b1_S1077 = 1077;
  localparam test_b1_S1078 = 1078;
  localparam test_b1_S1079 = 1079;
  localparam test_b1_S1080 = 1080;
  localparam test_b1_S1081 = 1081;
  localparam test_b1_S1082 = 1082;
  localparam test_b1_S1083 = 1083;
  localparam test_b1_S1084 = 1084;
  localparam test_b1_S1085 = 1085;
  localparam test_b1_S1086 = 1086;
  localparam test_b1_S1087 = 1087;
  localparam test_b1_S1088 = 1088;
  localparam test_b1_S1089 = 1089;
  localparam test_b1_S1090 = 1090;
  localparam test_b1_S1091 = 1091;
  localparam test_b1_S1092 = 1092;
  localparam test_b1_S1093 = 1093;
  localparam test_b1_S1094 = 1094;
  localparam test_b1_S1095 = 1095;
  localparam test_b1_S1096 = 1096;
  localparam test_b1_S1097 = 1097;
  localparam test_b1_S1098 = 1098;
  localparam test_b1_S1099 = 1099;
  localparam test_b1_S1100 = 1100;
  localparam test_b1_S1101 = 1101;
  localparam test_b1_S1102 = 1102;
  localparam test_b1_S1103 = 1103;
  localparam test_b1_S1104 = 1104;
  localparam test_b1_S1105 = 1105;
  localparam test_b1_S1106 = 1106;
  localparam test_b1_S1107 = 1107;
  localparam test_b1_S1108 = 1108;
  localparam test_b1_S1109 = 1109;
  localparam test_b1_S1110 = 1110;
  localparam test_b1_S1111 = 1111;
  localparam test_b1_S1112 = 1112;
  localparam test_b1_S1113 = 1113;
  localparam test_b1_S1114 = 1114;
  localparam test_b1_S1115 = 1115;
  localparam test_b1_S1116 = 1116;
  localparam test_b1_S1117 = 1117;
  localparam test_b1_S1118 = 1118;
  localparam test_b1_S1119 = 1119;
  localparam test_b1_S1120 = 1120;
  localparam test_b1_S1121 = 1121;
  localparam test_b1_S1122 = 1122;
  localparam test_b1_S1123 = 1123;
  localparam test_b1_S1124 = 1124;
  localparam test_b1_S1125 = 1125;
  localparam test_b1_S1126 = 1126;
  localparam test_b1_S1127 = 1127;
  localparam test_b1_S1128 = 1128;
  localparam test_b1_S1129 = 1129;
  localparam test_b1_S1130 = 1130;
  localparam test_b1_S1131 = 1131;
  localparam test_b1_S1132 = 1132;
  localparam test_b1_S1133 = 1133;
  localparam test_b1_S1134 = 1134;
  localparam test_b1_S1135 = 1135;
  localparam test_b1_S1136 = 1136;
  localparam test_b1_S1137 = 1137;
  localparam test_b1_S1138 = 1138;
  localparam test_b1_S1139 = 1139;
  localparam test_b1_S1140 = 1140;
  localparam test_b1_S1141 = 1141;
  localparam test_b1_S1142 = 1142;
  localparam test_b1_S1143 = 1143;
  localparam test_b1_S1144 = 1144;
  localparam test_b1_S1145 = 1145;
  localparam test_b1_S1146 = 1146;
  localparam test_b1_S1147 = 1147;
  localparam test_b1_S1148 = 1148;
  localparam test_b1_S1149 = 1149;
  localparam test_b1_S1150 = 1150;
  localparam test_b1_S1151 = 1151;
  localparam test_b1_S1152 = 1152;
  localparam test_b1_S1153 = 1153;
  localparam test_b1_S1154 = 1154;
  localparam test_b1_S1155 = 1155;
  localparam test_b1_S1156 = 1156;
  localparam test_b1_S1157 = 1157;
  localparam test_b1_S1158 = 1158;
  localparam test_b1_S1159 = 1159;
  localparam test_b1_S1160 = 1160;
  localparam test_b1_S1161 = 1161;
  localparam test_b1_S1162 = 1162;
  localparam test_b1_S1163 = 1163;
  localparam test_b1_S1164 = 1164;
  localparam test_b1_S1165 = 1165;
  localparam test_b1_S1166 = 1166;
  localparam test_b1_S1167 = 1167;
  localparam test_b1_S1168 = 1168;
  localparam test_b1_S1169 = 1169;
  localparam test_b1_S1170 = 1170;
  localparam test_b1_S1171 = 1171;
  localparam test_b1_S1172 = 1172;
  localparam test_b1_S1173 = 1173;
  localparam test_b1_S1174 = 1174;
  localparam test_b1_S1175 = 1175;
  localparam test_b1_S1176 = 1176;
  localparam test_b1_S1177 = 1177;
  localparam test_b1_S1178 = 1178;
  localparam test_b1_S1179 = 1179;
  localparam test_b1_S1180 = 1180;
  localparam test_b1_S1181 = 1181;
  localparam test_b1_S1182 = 1182;
  localparam test_b1_S1183 = 1183;
  localparam test_b1_S1184 = 1184;
  localparam test_b1_S1185 = 1185;
  localparam test_b1_S1186 = 1186;
  localparam test_b1_S1187 = 1187;
  localparam test_b1_S1188 = 1188;
  localparam test_b1_S1189 = 1189;
  localparam test_b1_S1190 = 1190;
  localparam test_b1_S1191 = 1191;
  localparam test_b1_S1192 = 1192;
  localparam test_b1_S1193 = 1193;
  localparam test_b1_S1194 = 1194;
  localparam test_b1_S1195 = 1195;
  localparam test_b1_S1196 = 1196;
  localparam test_b1_S1197 = 1197;
  localparam test_b1_S1198 = 1198;
  localparam test_b1_S1199 = 1199;
  localparam test_b1_S1200 = 1200;
  localparam test_b1_S1201 = 1201;
  localparam test_b1_S1202 = 1202;
  localparam test_b1_S1203 = 1203;
  localparam test_b1_S1204 = 1204;
  localparam test_b1_S1205 = 1205;
  localparam test_b1_S1206 = 1206;
  localparam test_b1_S1207 = 1207;
  localparam test_b1_S1208 = 1208;
  localparam test_b1_S1209 = 1209;
  localparam test_b1_S1210 = 1210;
  localparam test_b1_S1211 = 1211;
  localparam test_b1_S1212 = 1212;
  localparam test_b1_S1213 = 1213;
  localparam test_b1_S1214 = 1214;
  localparam test_b1_S1215 = 1215;
  localparam test_b1_S1216 = 1216;
  localparam test_b1_S1217 = 1217;
  localparam test_b1_S1218 = 1218;
  localparam test_b1_S1219 = 1219;
  localparam test_b1_S1220 = 1220;
  localparam test_b1_S1221 = 1221;
  localparam test_b1_S1222 = 1222;
  localparam test_b1_S1223 = 1223;
  localparam test_b1_S1224 = 1224;
  localparam test_b1_S1225 = 1225;
  localparam test_b1_S1226 = 1226;
  localparam test_b1_S1227 = 1227;
  localparam test_b1_S1228 = 1228;
  localparam test_b1_S1229 = 1229;
  localparam test_b1_S1230 = 1230;
  localparam test_b1_S1231 = 1231;
  localparam test_b1_S1232 = 1232;
  localparam test_b1_S1233 = 1233;
  localparam test_b1_S1234 = 1234;
  localparam test_b1_S1235 = 1235;
  localparam test_b1_S1236 = 1236;
  localparam test_b1_S1237 = 1237;
  localparam test_b1_S1238 = 1238;
  localparam test_b1_S1239 = 1239;
  localparam test_b1_S1240 = 1240;
  localparam test_b1_S1241 = 1241;
  localparam test_b1_S1242 = 1242;
  localparam test_b1_S1243 = 1243;
  localparam test_b1_S1244 = 1244;
  localparam test_b1_S1245 = 1245;
  localparam test_b1_S1246 = 1246;
  localparam test_b1_S1247 = 1247;
  localparam test_b1_S1248 = 1248;
  localparam test_b1_S1249 = 1249;
  localparam test_b1_S1250 = 1250;
  localparam test_b1_S1251 = 1251;
  localparam test_b1_S1252 = 1252;
  localparam test_b1_S1253 = 1253;
  localparam test_b1_S1254 = 1254;
  localparam test_b1_S1255 = 1255;
  localparam test_b1_S1256 = 1256;
  localparam test_b1_S1257 = 1257;
  localparam test_b1_S1258 = 1258;
  localparam test_b1_S1259 = 1259;
  localparam test_b1_S1260 = 1260;
  localparam test_b1_S1261 = 1261;
  localparam test_b1_S1262 = 1262;
  localparam test_b1_S1263 = 1263;
  localparam test_b1_S1264 = 1264;
  localparam test_b1_S1265 = 1265;
  localparam test_b1_S1266 = 1266;
  localparam test_b1_S1267 = 1267;
  localparam test_b1_S1268 = 1268;
  localparam test_b1_S1269 = 1269;
  localparam test_b1_S1270 = 1270;
  localparam test_b1_S1271 = 1271;
  localparam test_b1_S1272 = 1272;
  localparam test_b1_S1273 = 1273;
  localparam test_b1_S1274 = 1274;
  localparam test_b1_S1275 = 1275;
  localparam test_b1_S1276 = 1276;
  localparam test_b1_S1277 = 1277;
  localparam test_b1_S1278 = 1278;
  localparam test_b1_S1279 = 1279;
  localparam test_b1_S1280 = 1280;
  localparam test_b1_S1281 = 1281;
  localparam test_b1_S1282 = 1282;
  localparam test_b1_S1283 = 1283;
  localparam test_b1_S1284 = 1284;
  localparam test_b1_S1285 = 1285;
  localparam test_b1_S1286 = 1286;
  localparam test_b1_S1287 = 1287;
  localparam test_b1_S1288 = 1288;
  localparam test_b1_S1289 = 1289;
  localparam test_b1_S1290 = 1290;
  localparam test_b1_S1291 = 1291;
  localparam test_b1_S1292 = 1292;
  localparam test_b1_S1293 = 1293;
  localparam test_b1_S1294 = 1294;
  localparam test_b1_S1295 = 1295;
  localparam test_b1_S1296 = 1296;
  localparam test_b1_S1297 = 1297;
  localparam test_b1_S1298 = 1298;
  localparam test_b1_S1299 = 1299;
  localparam test_b1_S1300 = 1300;
  localparam test_b1_S1301 = 1301;
  localparam test_b1_S1302 = 1302;
  localparam test_b1_S1303 = 1303;
  localparam test_b1_S1304 = 1304;
  localparam test_b1_S1305 = 1305;
  localparam test_b1_S1306 = 1306;
  localparam test_b1_S1307 = 1307;
  localparam test_b1_S1308 = 1308;
  localparam test_b1_S1309 = 1309;
  localparam test_b1_S1310 = 1310;
  localparam test_b1_S1311 = 1311;
  localparam test_b1_S1312 = 1312;
  localparam test_b1_S1313 = 1313;
  localparam test_b1_S1314 = 1314;
  localparam test_b1_S1315 = 1315;
  localparam test_b1_S1316 = 1316;
  localparam test_b1_S1317 = 1317;
  localparam test_b1_S1318 = 1318;
  localparam test_b1_S1319 = 1319;
  localparam test_b1_S1320 = 1320;
  localparam test_b1_S1321 = 1321;
  localparam test_b1_S1322 = 1322;
  localparam test_b1_S1323 = 1323;
  localparam test_b1_S1324 = 1324;
  localparam test_b1_S1325 = 1325;
  localparam test_b1_S1326 = 1326;
  localparam test_b1_S1327 = 1327;
  localparam test_b1_S1328 = 1328;
  localparam test_b1_S1329 = 1329;
  localparam test_b1_S1330 = 1330;
  localparam test_b1_S1331 = 1331;
  localparam test_b1_S1332 = 1332;
  localparam test_b1_S1333 = 1333;
  localparam test_b1_S1334 = 1334;
  localparam test_b1_S1335 = 1335;
  localparam test_b1_S1336 = 1336;
  localparam test_b1_S1337 = 1337;
  localparam test_b1_S1338 = 1338;
  localparam test_b1_S1339 = 1339;
  localparam test_b1_S1340 = 1340;
  localparam test_b1_S1341 = 1341;
  localparam test_b1_S1342 = 1342;
  localparam test_b1_S1343 = 1343;
  localparam test_b1_S1344 = 1344;
  localparam test_b1_S1345 = 1345;
  localparam test_b1_S1346 = 1346;
  localparam test_b1_S1347 = 1347;
  localparam test_b1_S1348 = 1348;
  localparam test_b1_S1349 = 1349;
  localparam test_b1_S1350 = 1350;
  localparam test_b1_S1351 = 1351;
  localparam test_b1_S1352 = 1352;
  localparam test_b1_S1353 = 1353;
  localparam test_b1_S1354 = 1354;
  localparam test_b1_S1355 = 1355;
  localparam test_b1_S1356 = 1356;
  localparam test_b1_S1357 = 1357;
  localparam test_b1_S1358 = 1358;
  localparam test_b1_S1359 = 1359;
  localparam test_b1_S1360 = 1360;
  localparam test_b1_S1361 = 1361;
  localparam test_b1_S1362 = 1362;
  localparam test_b1_S1363 = 1363;
  localparam test_b1_S1364 = 1364;
  localparam test_b1_S1365 = 1365;
  localparam test_b1_S1366 = 1366;
  localparam test_b1_S1367 = 1367;
  localparam test_b1_S1368 = 1368;
  localparam test_b1_S1369 = 1369;
  localparam test_b1_S1370 = 1370;
  localparam test_b1_S1371 = 1371;
  localparam test_b1_S1372 = 1372;
  localparam test_b1_S1373 = 1373;
  localparam test_b1_S1374 = 1374;
  localparam test_b1_S1375 = 1375;
  localparam test_b1_S1376 = 1376;
  localparam test_b1_S1377 = 1377;
  localparam test_b1_S1378 = 1378;
  localparam test_b1_S1379 = 1379;
  localparam test_b1_S1380 = 1380;
  localparam test_b1_S1381 = 1381;
  localparam test_b1_S1382 = 1382;
  localparam test_b1_S1383 = 1383;
  localparam test_b1_S1384 = 1384;
  localparam test_b1_S1385 = 1385;
  localparam test_b1_S1386 = 1386;
  localparam test_b1_S1387 = 1387;
  localparam test_b1_S1388 = 1388;
  localparam test_b1_S1389 = 1389;
  localparam test_b1_S1390 = 1390;
  localparam test_b1_S1391 = 1391;
  localparam test_b1_S1392 = 1392;
  localparam test_b1_S1393 = 1393;
  localparam test_b1_S1394 = 1394;
  localparam test_b1_S1395 = 1395;
  localparam test_b1_S1396 = 1396;
  localparam test_b1_S1397 = 1397;
  localparam test_b1_S1398 = 1398;
  localparam test_b1_S1399 = 1399;
  localparam test_b1_S1400 = 1400;
  localparam test_b1_S1401 = 1401;
  localparam test_b1_S1402 = 1402;
  localparam test_b1_S1403 = 1403;
  localparam test_b1_S1404 = 1404;
  localparam test_b1_S1405 = 1405;
  localparam test_b1_S1406 = 1406;
  localparam test_b1_S1407 = 1407;
  localparam test_b1_S1408 = 1408;
  localparam test_b1_S1409 = 1409;
  localparam test_b1_S1410 = 1410;
  localparam test_b1_S1411 = 1411;
  localparam test_b1_S1412 = 1412;
  localparam test_b1_S1413 = 1413;
  localparam test_b1_S1414 = 1414;
  localparam test_b1_S1415 = 1415;
  localparam test_b1_S1416 = 1416;
  localparam test_b1_S1417 = 1417;
  localparam test_b1_S1418 = 1418;
  localparam test_b1_S1419 = 1419;
  localparam test_b1_S1420 = 1420;
  localparam test_b1_S1421 = 1421;
  localparam test_b1_S1422 = 1422;
  localparam test_b1_S1423 = 1423;
  localparam test_b1_S1424 = 1424;
  localparam test_b1_S1425 = 1425;
  localparam test_b1_S1426 = 1426;
  localparam test_b1_S1427 = 1427;
  localparam test_b1_S1428 = 1428;
  localparam test_b1_S1429 = 1429;
  localparam test_b1_S1430 = 1430;
  localparam test_b1_S1431 = 1431;
  localparam test_b1_S1432 = 1432;
  localparam test_b1_S1433 = 1433;
  localparam test_b1_S1434 = 1434;
  localparam test_b1_S1435 = 1435;
  localparam test_b1_S1436 = 1436;
  localparam test_b1_S1437 = 1437;
  localparam test_b1_S1438 = 1438;
  localparam test_b1_S1439 = 1439;
  localparam test_b1_S1440 = 1440;
  localparam test_b1_S1441 = 1441;
  localparam test_b1_S1442 = 1442;
  localparam test_b1_S1443 = 1443;
  localparam test_b1_S1444 = 1444;
  localparam test_b1_S1445 = 1445;
  localparam test_b1_S1446 = 1446;
  localparam test_b1_S1447 = 1447;
  localparam test_b1_S1448 = 1448;
  localparam test_b1_S1449 = 1449;
  localparam test_b1_S1450 = 1450;
  localparam test_b1_S1451 = 1451;
  localparam test_b1_S1452 = 1452;
  localparam test_b1_S1453 = 1453;
  localparam test_b1_S1454 = 1454;
  localparam test_b1_S1455 = 1455;
  localparam test_b1_S1456 = 1456;
  localparam test_b1_S1457 = 1457;
  localparam test_b1_S1458 = 1458;
  localparam test_b1_S1459 = 1459;
  localparam test_b1_S1460 = 1460;
  localparam test_b1_S1461 = 1461;
  localparam test_b1_S1462 = 1462;
  localparam test_b1_S1463 = 1463;
  localparam test_b1_S1464 = 1464;
  localparam test_b1_S1465 = 1465;
  localparam test_b1_S1466 = 1466;
  localparam test_b1_S1467 = 1467;
  localparam test_b1_S1468 = 1468;
  localparam test_b1_S1469 = 1469;
  localparam test_b1_S1470 = 1470;
  localparam test_b1_S1471 = 1471;
  localparam test_b1_S1472 = 1472;
  localparam test_b1_S1473 = 1473;
  localparam test_b1_S1474 = 1474;
  localparam test_b1_S1475 = 1475;
  localparam test_b1_S1476 = 1476;
  localparam test_b1_S1477 = 1477;
  localparam test_b1_S1478 = 1478;
  localparam test_b1_S1479 = 1479;
  localparam test_b1_S1480 = 1480;
  localparam test_b1_S1481 = 1481;
  localparam test_b1_S1482 = 1482;
  localparam test_b1_S1483 = 1483;
  localparam test_b1_S1484 = 1484;
  localparam test_b1_S1485 = 1485;
  localparam test_b1_S1486 = 1486;
  localparam test_b1_S1487 = 1487;
  localparam test_b1_S1488 = 1488;
  localparam test_b1_S1489 = 1489;
  localparam test_b1_S1490 = 1490;
  localparam test_b1_S1491 = 1491;
  localparam test_b1_S1492 = 1492;
  localparam test_b1_S1493 = 1493;
  localparam test_b1_S1494 = 1494;
  localparam test_b1_S1495 = 1495;
  localparam test_b1_S1496 = 1496;
  localparam test_b1_S1497 = 1497;
  localparam test_b1_S1498 = 1498;
  localparam test_b1_S1499 = 1499;
  localparam test_b1_S1500 = 1500;
  localparam test_b1_S1501 = 1501;
  localparam test_b1_S1502 = 1502;
  localparam test_b1_S1503 = 1503;
  localparam test_b1_S1504 = 1504;
  localparam test_b1_S1505 = 1505;
  localparam test_b1_S1506 = 1506;
  localparam test_b1_S1507 = 1507;
  localparam test_b1_S1508 = 1508;
  localparam test_b1_S1509 = 1509;
  localparam test_b1_S1510 = 1510;
  localparam test_b1_S1511 = 1511;
  localparam test_b1_S1512 = 1512;
  localparam test_b1_S1513 = 1513;
  localparam test_b1_S1514 = 1514;
  localparam test_b1_S1515 = 1515;
  localparam test_b1_S1516 = 1516;
  localparam test_b1_S1517 = 1517;
  localparam test_b1_S1518 = 1518;
  localparam test_b1_S1519 = 1519;
  localparam test_b1_S1520 = 1520;
  localparam test_b1_S1521 = 1521;
  localparam test_b1_S1522 = 1522;
  localparam test_b1_S1523 = 1523;
  localparam test_b1_S1524 = 1524;
  localparam test_b1_S1525 = 1525;
  localparam test_b1_S1526 = 1526;
  localparam test_b1_S1527 = 1527;
  localparam test_b1_S1528 = 1528;
  localparam test_b1_S1529 = 1529;
  localparam test_b1_S1530 = 1530;
  localparam test_b1_S1531 = 1531;
  localparam test_b1_S1532 = 1532;
  localparam test_b1_S1533 = 1533;
  localparam test_b1_S1534 = 1534;
  localparam test_b1_S1535 = 1535;
  localparam test_b1_S1536 = 1536;
  localparam test_b1_S1537 = 1537;
  localparam test_b1_S1538 = 1538;
  localparam test_b1_S1539 = 1539;
  localparam test_b1_S1540 = 1540;
  localparam test_b1_S1541 = 1541;
  localparam test_b1_S1542 = 1542;
  localparam test_b1_S1543 = 1543;
  localparam test_b1_S1544 = 1544;
  localparam test_b1_S1545 = 1545;
  localparam test_b1_S1546 = 1546;
  localparam test_b1_S1547 = 1547;
  localparam test_b1_S1548 = 1548;
  localparam test_b1_S1549 = 1549;
  localparam test_b1_S1550 = 1550;
  localparam test_b1_S1551 = 1551;
  localparam test_b1_S1552 = 1552;
  localparam test_b1_S1553 = 1553;
  localparam test_b1_S1554 = 1554;
  localparam test_b1_S1555 = 1555;
  localparam test_b1_S1556 = 1556;
  localparam test_b1_S1557 = 1557;
  localparam test_b1_S1558 = 1558;
  localparam test_b1_S1559 = 1559;
  localparam test_b1_S1560 = 1560;
  localparam test_b1_S1561 = 1561;
  localparam test_b1_S1562 = 1562;
  localparam test_b1_S1563 = 1563;
  localparam test_b1_S1564 = 1564;
  localparam test_b1_S1565 = 1565;
  localparam test_b1_S1566 = 1566;
  localparam test_b1_S1567 = 1567;
  localparam test_b1_S1568 = 1568;
  localparam test_b1_S1569 = 1569;
  localparam test_b1_S1570 = 1570;
  localparam test_b1_S1571 = 1571;
  localparam test_b1_S1572 = 1572;
  localparam test_b1_S1573 = 1573;
  localparam test_b1_S1574 = 1574;
  localparam test_b1_S1575 = 1575;
  localparam test_b1_S1576 = 1576;
  localparam test_b1_S1577 = 1577;
  localparam test_b1_S1578 = 1578;
  localparam test_b1_S1579 = 1579;
  localparam test_b1_S1580 = 1580;
  localparam test_b1_S1581 = 1581;
  localparam test_b1_S1582 = 1582;
  localparam test_b1_S1583 = 1583;
  localparam test_b1_S1584 = 1584;
  localparam test_b1_S1585 = 1585;
  localparam test_b1_S1586 = 1586;
  localparam test_b1_S1587 = 1587;
  localparam test_b1_S1588 = 1588;
  localparam test_b1_S1589 = 1589;
  localparam test_b1_S1590 = 1590;
  localparam test_b1_S1591 = 1591;
  localparam test_b1_S1592 = 1592;
  localparam test_b1_S1593 = 1593;
  localparam test_b1_S1594 = 1594;
  localparam test_b1_S1595 = 1595;
  localparam test_b1_S1596 = 1596;
  localparam test_b1_S1597 = 1597;
  localparam test_b1_S1598 = 1598;
  localparam test_b1_S1599 = 1599;
  localparam test_b1_S1600 = 1600;
  localparam test_b1_S1601 = 1601;
  localparam test_b1_S1602 = 1602;
  localparam test_b1_S1603 = 1603;
  localparam test_b1_S1604 = 1604;
  localparam test_b1_S1605 = 1605;
  localparam test_b1_S1606 = 1606;
  localparam test_b1_S1607 = 1607;
  localparam test_b1_S1608 = 1608;
  localparam test_b1_S1609 = 1609;
  localparam test_b1_S1610 = 1610;
  localparam test_b1_S1611 = 1611;
  localparam test_b1_S1612 = 1612;
  localparam test_b1_S1613 = 1613;
  localparam test_b1_S1614 = 1614;
  localparam test_b1_S1615 = 1615;
  localparam test_b1_S1616 = 1616;
  localparam test_b1_S1617 = 1617;
  localparam test_b1_S1618 = 1618;
  localparam test_b1_S1619 = 1619;
  localparam test_b1_S1620 = 1620;
  localparam test_b1_S1621 = 1621;
  localparam test_b1_S1622 = 1622;
  localparam test_b1_S1623 = 1623;
  localparam test_b1_S1624 = 1624;
  localparam test_b1_S1625 = 1625;
  localparam test_b1_S1626 = 1626;
  localparam test_b1_S1627 = 1627;
  localparam test_b1_S1628 = 1628;
  localparam test_b1_S1629 = 1629;
  localparam test_b1_S1630 = 1630;
  localparam test_b1_S1631 = 1631;
  localparam test_b1_S1632 = 1632;
  localparam test_b1_S1633 = 1633;
  localparam test_b1_S1634 = 1634;
  localparam test_b1_S1635 = 1635;
  localparam test_b1_S1636 = 1636;
  localparam test_b1_S1637 = 1637;
  localparam test_b1_S1638 = 1638;
  localparam test_b1_S1639 = 1639;
  localparam test_b1_S1640 = 1640;
  localparam test_b1_S1641 = 1641;
  localparam test_b1_S1642 = 1642;
  localparam test_b1_S1643 = 1643;
  localparam test_b1_S1644 = 1644;
  localparam test_b1_S1645 = 1645;
  localparam test_b1_S1646 = 1646;
  localparam test_b1_S1647 = 1647;
  localparam test_b1_S1648 = 1648;
  localparam test_b1_S1649 = 1649;
  localparam test_b1_S1650 = 1650;
  localparam test_b1_S1651 = 1651;
  localparam test_b1_S1652 = 1652;
  localparam test_b1_S1653 = 1653;
  localparam test_b1_S1654 = 1654;
  localparam test_b1_S1655 = 1655;
  localparam test_b1_S1656 = 1656;
  localparam test_b1_S1657 = 1657;
  localparam test_b1_S1658 = 1658;
  localparam test_b1_S1659 = 1659;
  localparam test_b1_S1660 = 1660;
  localparam test_b1_S1661 = 1661;
  localparam test_b1_S1662 = 1662;
  localparam test_b1_S1663 = 1663;
  localparam test_b1_S1664 = 1664;
  localparam test_b1_S1665 = 1665;
  localparam test_b1_S1666 = 1666;
  localparam test_b1_S1667 = 1667;
  localparam test_b1_S1668 = 1668;
  localparam test_b1_S1669 = 1669;
  localparam test_b1_S1670 = 1670;
  localparam test_b1_S1671 = 1671;
  localparam test_b1_S1672 = 1672;
  localparam test_b1_S1673 = 1673;
  localparam test_b1_S1674 = 1674;
  localparam test_b1_S1675 = 1675;
  localparam test_b1_S1676 = 1676;
  localparam test_b1_S1677 = 1677;
  localparam test_b1_S1678 = 1678;
  localparam test_b1_S1679 = 1679;
  localparam test_b1_S1680 = 1680;
  localparam test_b1_S1681 = 1681;
  localparam test_b1_S1682 = 1682;
  localparam test_b1_S1683 = 1683;
  localparam test_b1_S1684 = 1684;
  localparam test_b1_S1685 = 1685;
  localparam test_b1_S1686 = 1686;
  localparam test_b1_S1687 = 1687;
  localparam test_b1_S1688 = 1688;
  localparam test_b1_S1689 = 1689;
  localparam test_b1_S1690 = 1690;
  localparam test_b1_S1691 = 1691;
  localparam test_b1_S1692 = 1692;
  localparam test_b1_S1693 = 1693;
  localparam test_b1_S1694 = 1694;
  localparam test_b1_S1695 = 1695;
  localparam test_b1_S1696 = 1696;
  localparam test_b1_S1697 = 1697;
  localparam test_b1_S1698 = 1698;
  localparam test_b1_S1699 = 1699;
  localparam test_b1_S1700 = 1700;
  localparam test_b1_S1701 = 1701;
  localparam test_b1_S1702 = 1702;
  localparam test_b1_S1703 = 1703;
  localparam test_b1_S1704 = 1704;
  localparam test_b1_S1705 = 1705;
  localparam test_b1_S1706 = 1706;
  localparam test_b1_S1707 = 1707;
  localparam test_b1_S1708 = 1708;
  localparam test_b1_S1709 = 1709;
  localparam test_b1_S1710 = 1710;
  localparam test_b1_S1711 = 1711;
  localparam test_b1_S1712 = 1712;
  localparam test_b1_S1713 = 1713;
  localparam test_b1_S1714 = 1714;
  localparam test_b1_S1715 = 1715;
  localparam test_b1_S1716 = 1716;
  localparam test_b1_S1717 = 1717;
  localparam test_b1_S1718 = 1718;
  localparam test_b1_S1719 = 1719;
  localparam test_b1_S1720 = 1720;
  localparam test_b1_S1721 = 1721;
  localparam test_b1_S1722 = 1722;
  localparam test_b1_S1723 = 1723;
  localparam test_b1_S1724 = 1724;
  localparam test_b1_S1725 = 1725;
  localparam test_b1_S1726 = 1726;
  localparam test_b1_S1727 = 1727;
  localparam test_b1_S1728 = 1728;
  localparam test_b1_S1729 = 1729;
  localparam test_b1_S1730 = 1730;
  localparam test_b1_S1731 = 1731;
  localparam test_b1_S1732 = 1732;
  localparam test_b1_S1733 = 1733;
  localparam test_b1_S1734 = 1734;
  localparam test_b1_S1735 = 1735;
  localparam test_b1_S1736 = 1736;
  localparam test_b1_S1737 = 1737;
  localparam test_b1_S1738 = 1738;
  localparam test_b1_S1739 = 1739;
  localparam test_b1_S1740 = 1740;
  localparam test_b1_S1741 = 1741;
  localparam test_b1_S1742 = 1742;
  localparam test_b1_S1743 = 1743;
  localparam test_b1_S1744 = 1744;
  localparam test_b1_S1745 = 1745;
  localparam test_b1_S1746 = 1746;
  localparam test_b1_S1747 = 1747;
  localparam test_b1_S1748 = 1748;
  localparam test_b1_S1749 = 1749;
  localparam test_b1_S1750 = 1750;
  localparam test_b1_S1751 = 1751;
  localparam test_b1_S1752 = 1752;
  localparam test_b1_S1753 = 1753;
  localparam test_b1_S1754 = 1754;
  localparam test_b1_S1755 = 1755;
  localparam test_b1_S1756 = 1756;
  localparam test_b1_S1757 = 1757;
  localparam test_b1_S1758 = 1758;
  localparam test_b1_S1759 = 1759;
  localparam test_b1_S1760 = 1760;
  localparam test_b1_S1761 = 1761;
  localparam test_b1_S1762 = 1762;
  localparam test_b1_S1763 = 1763;
  localparam test_b1_S1764 = 1764;
  localparam test_b1_S1765 = 1765;
  localparam test_b1_S1766 = 1766;
  localparam test_b1_S1767 = 1767;
  localparam test_b1_S1768 = 1768;
  localparam test_b1_S1769 = 1769;
  localparam test_b1_S1770 = 1770;
  localparam test_b1_S1771 = 1771;
  localparam test_b1_S1772 = 1772;
  localparam test_b1_S1773 = 1773;
  localparam test_b1_S1774 = 1774;
  localparam test_b1_S1775 = 1775;
  localparam test_b1_S1776 = 1776;
  localparam test_b1_S1777 = 1777;
  localparam test_b1_S1778 = 1778;
  localparam test_b1_S1779 = 1779;
  localparam test_b1_S1780 = 1780;
  localparam test_b1_S1781 = 1781;
  localparam test_b1_S1782 = 1782;
  localparam test_b1_S1783 = 1783;
  localparam test_b1_S1784 = 1784;
  localparam test_b1_S1785 = 1785;
  localparam test_b1_S1786 = 1786;
  localparam test_b1_S1787 = 1787;
  localparam test_b1_S1788 = 1788;
  localparam test_b1_S1789 = 1789;
  localparam test_b1_S1790 = 1790;
  localparam test_b1_S1791 = 1791;
  localparam test_b1_S1792 = 1792;
  localparam test_b1_S1793 = 1793;
  localparam test_b1_S1794 = 1794;
  localparam test_b1_S1795 = 1795;
  localparam test_b1_S1796 = 1796;
  localparam test_b1_S1797 = 1797;
  localparam test_b1_S1798 = 1798;
  localparam test_b1_S1799 = 1799;
  localparam test_b1_S1800 = 1800;
  localparam test_b1_S1801 = 1801;
  localparam test_b1_S1802 = 1802;
  localparam test_b1_S1803 = 1803;
  localparam test_b1_S1804 = 1804;
  localparam test_b1_S1805 = 1805;
  localparam test_b1_S1806 = 1806;
  localparam test_b1_S1807 = 1807;
  localparam test_b1_S1808 = 1808;
  localparam test_b1_S1809 = 1809;
  localparam test_b1_S1810 = 1810;
  localparam test_b1_S1811 = 1811;
  localparam test_b1_S1812 = 1812;
  localparam test_b1_S1813 = 1813;
  localparam test_b1_S1814 = 1814;
  localparam test_b1_S1815 = 1815;
  localparam test_b1_S1816 = 1816;
  localparam test_b1_S1817 = 1817;
  localparam test_b1_S1818 = 1818;
  localparam test_b1_S1819 = 1819;
  localparam test_b1_S1820 = 1820;
  localparam test_b1_S1821 = 1821;
  localparam test_b1_S1822 = 1822;
  localparam test_b1_S1823 = 1823;
  localparam test_b1_S1824 = 1824;
  localparam test_b1_S1825 = 1825;
  localparam test_b1_S1826 = 1826;
  localparam test_b1_S1827 = 1827;
  localparam test_b1_S1828 = 1828;
  localparam test_b1_S1829 = 1829;
  localparam test_b1_S1830 = 1830;
  localparam test_b1_S1831 = 1831;
  localparam test_b1_S1832 = 1832;
  localparam test_b1_S1833 = 1833;
  localparam test_b1_S1834 = 1834;
  localparam test_b1_S1835 = 1835;
  localparam test_b1_S1836 = 1836;
  localparam test_b1_S1837 = 1837;
  localparam test_b1_S1838 = 1838;
  localparam test_b1_S1839 = 1839;
  localparam test_b1_S1840 = 1840;
  localparam test_b1_S1841 = 1841;
  localparam test_b1_S1842 = 1842;
  localparam test_b1_S1843 = 1843;
  localparam test_b1_S1844 = 1844;
  localparam test_b1_S1845 = 1845;
  localparam test_b1_S1846 = 1846;
  localparam test_b1_S1847 = 1847;
  localparam test_b1_S1848 = 1848;
  localparam test_b1_S1849 = 1849;
  localparam test_b1_S1850 = 1850;
  localparam test_b1_S1851 = 1851;
  localparam test_b1_S1852 = 1852;
  localparam test_b1_S1853 = 1853;
  localparam test_b1_S1854 = 1854;
  localparam test_b1_S1855 = 1855;
  localparam test_b1_S1856 = 1856;
  localparam test_b1_S1857 = 1857;
  localparam test_b1_S1858 = 1858;
  localparam test_b1_S1859 = 1859;
  localparam test_b1_S1860 = 1860;
  localparam test_b1_S1861 = 1861;
  localparam test_b1_S1862 = 1862;
  localparam test_b1_S1863 = 1863;
  localparam test_b1_S1864 = 1864;
  localparam test_b1_S1865 = 1865;
  localparam test_b1_S1866 = 1866;
  localparam test_b1_S1867 = 1867;
  localparam test_b1_S1868 = 1868;
  localparam test_b1_S1869 = 1869;
  localparam test_b1_S1870 = 1870;
  localparam test_b1_S1871 = 1871;
  localparam test_b1_S1872 = 1872;
  localparam test_b1_S1873 = 1873;
  localparam test_b1_S1874 = 1874;
  localparam test_b1_S1875 = 1875;
  localparam test_b1_S1876 = 1876;
  localparam test_b1_S1877 = 1877;
  localparam test_b1_S1878 = 1878;
  localparam test_b1_S1879 = 1879;
  localparam test_b1_S1880 = 1880;
  localparam test_b1_S1881 = 1881;
  localparam test_b1_S1882 = 1882;
  localparam test_b1_S1883 = 1883;
  localparam test_b1_S1884 = 1884;
  localparam test_b1_S1885 = 1885;
  localparam test_b1_S1886 = 1886;
  localparam test_b1_S1887 = 1887;
  localparam test_b1_S1888 = 1888;
  localparam test_b1_S1889 = 1889;
  localparam test_b1_S1890 = 1890;
  localparam test_b1_S1891 = 1891;
  localparam test_b1_S1892 = 1892;
  localparam test_b1_S1893 = 1893;
  localparam test_b1_S1894 = 1894;
  localparam test_b1_S1895 = 1895;
  localparam test_b1_S1896 = 1896;
  localparam test_b1_S1897 = 1897;
  localparam test_b1_S1898 = 1898;
  localparam test_b1_S1899 = 1899;
  localparam test_b1_S1900 = 1900;
  localparam test_b1_S1901 = 1901;
  localparam test_b1_S1902 = 1902;
  localparam test_b1_S1903 = 1903;
  localparam test_b1_S1904 = 1904;
  localparam test_b1_S1905 = 1905;
  localparam test_b1_S1906 = 1906;
  localparam test_b1_S1907 = 1907;
  localparam test_b1_S1908 = 1908;
  localparam test_b1_S1909 = 1909;
  localparam test_b1_S1910 = 1910;
  localparam test_b1_S1911 = 1911;
  localparam test_b1_S1912 = 1912;
  localparam test_b1_S1913 = 1913;
  localparam test_b1_S1914 = 1914;
  localparam test_b1_S1915 = 1915;
  localparam test_b1_S1916 = 1916;
  localparam test_b1_S1917 = 1917;
  localparam test_b1_S1918 = 1918;
  localparam test_b1_S1919 = 1919;
  localparam test_b1_S1920 = 1920;
  localparam test_b1_S1921 = 1921;
  localparam test_b1_S1922 = 1922;
  localparam test_b1_S1923 = 1923;
  localparam test_b1_S1924 = 1924;
  localparam test_b1_S1925 = 1925;
  localparam test_b1_S1926 = 1926;
  localparam test_b1_S1927 = 1927;
  localparam test_b1_S1928 = 1928;
  localparam test_b1_S1929 = 1929;
  localparam test_b1_S1930 = 1930;
  localparam test_b1_S1931 = 1931;
  localparam test_b1_S1932 = 1932;
  localparam test_b1_S1933 = 1933;
  localparam test_b1_S1934 = 1934;
  localparam test_b1_S1935 = 1935;
  localparam test_b1_S1936 = 1936;
  localparam test_b1_S1937 = 1937;
  localparam test_b1_S1938 = 1938;
  localparam test_b1_S1939 = 1939;
  localparam test_b1_S1940 = 1940;
  localparam test_b1_S1941 = 1941;
  localparam test_b1_S1942 = 1942;
  localparam test_b1_S1943 = 1943;
  localparam test_b1_S1944 = 1944;
  localparam test_b1_S1945 = 1945;
  localparam test_b1_S1946 = 1946;
  localparam test_b1_S1947 = 1947;
  localparam test_b1_S1948 = 1948;
  localparam test_b1_S1949 = 1949;
  localparam test_b1_S1950 = 1950;
  localparam test_b1_S1951 = 1951;
  localparam test_b1_S1952 = 1952;
  localparam test_b1_S1953 = 1953;
  localparam test_b1_S1954 = 1954;
  localparam test_b1_S1955 = 1955;
  localparam test_b1_S1956 = 1956;
  localparam test_b1_S1957 = 1957;
  localparam test_b1_S1958 = 1958;
  localparam test_b1_S1959 = 1959;
  localparam test_b1_S1960 = 1960;
  localparam test_b1_S1961 = 1961;
  localparam test_b1_S1962 = 1962;
  localparam test_b1_S1963 = 1963;
  localparam test_b1_S1964 = 1964;
  localparam test_b1_S1965 = 1965;
  localparam test_b1_S1966 = 1966;
  localparam test_b1_S1967 = 1967;
  localparam test_b1_S1968 = 1968;
  localparam test_b1_S1969 = 1969;
  localparam test_b1_S1970 = 1970;
  localparam test_b1_S1971 = 1971;
  localparam test_b1_S1972 = 1972;
  localparam test_b1_S1973 = 1973;
  localparam test_b1_S1974 = 1974;
  localparam test_b1_S1975 = 1975;
  localparam test_b1_S1976 = 1976;
  localparam test_b1_S1977 = 1977;
  localparam test_b1_S1978 = 1978;
  localparam test_b1_S1979 = 1979;
  localparam test_b1_S1980 = 1980;
  localparam test_b1_S1981 = 1981;
  localparam test_b1_S1982 = 1982;
  localparam test_b1_S1983 = 1983;
  localparam test_b1_S1984 = 1984;
  localparam test_b1_S1985 = 1985;
  localparam test_b1_S1986 = 1986;
  localparam test_b1_S1987 = 1987;
  localparam test_b1_S1988 = 1988;
  localparam test_b1_S1989 = 1989;
  localparam test_b1_S1990 = 1990;
  localparam test_b1_S1991 = 1991;
  localparam test_b1_S1992 = 1992;
  localparam test_b1_S1993 = 1993;
  localparam test_b1_S1994 = 1994;
  localparam test_b1_S1995 = 1995;
  localparam test_b1_S1996 = 1996;
  localparam test_b1_S1997 = 1997;
  localparam test_b1_S1998 = 1998;
  localparam test_b1_S1999 = 1999;
  localparam test_b1_S2000 = 2000;
  localparam test_b1_S2001 = 2001;
  localparam test_b1_S2002 = 2002;
  localparam test_b1_S2003 = 2003;
  localparam test_b1_S2004 = 2004;
  localparam test_b1_S2005 = 2005;
  localparam test_b1_S2006 = 2006;
  localparam test_b1_S2007 = 2007;
  localparam test_b1_S2008 = 2008;
  localparam test_b1_S2009 = 2009;
  localparam test_b1_S2010 = 2010;
  localparam test_b1_S2011 = 2011;
  localparam test_b1_S2012 = 2012;
  localparam test_b1_S2013 = 2013;
  localparam test_b1_S2014 = 2014;
  localparam test_b1_S2015 = 2015;
  localparam test_b1_S2016 = 2016;
  localparam test_b1_S2017 = 2017;
  localparam test_b1_S2018 = 2018;
  localparam test_b1_S2019 = 2019;
  localparam test_b1_S2020 = 2020;
  localparam test_b1_S2021 = 2021;
  localparam test_b1_S2022 = 2022;
  localparam test_b1_S2023 = 2023;
  localparam test_b1_S2024 = 2024;
  localparam test_b1_S2025 = 2025;
  localparam test_b1_S2026 = 2026;
  localparam test_b1_S2027 = 2027;
  localparam test_b1_S2028 = 2028;
  localparam test_b1_S2029 = 2029;
  localparam test_b1_S2030 = 2030;
  localparam test_b1_S2031 = 2031;
  localparam test_b1_S2032 = 2032;
  localparam test_b1_S2033 = 2033;
  localparam test_b1_S2034 = 2034;
  localparam test_b1_S2035 = 2035;
  localparam test_b1_S2036 = 2036;
  localparam test_b1_S2037 = 2037;
  localparam test_b1_S2038 = 2038;
  localparam test_b1_S2039 = 2039;
  localparam test_b1_S2040 = 2040;
  localparam test_b1_S2041 = 2041;
  localparam test_b1_S2042 = 2042;
  localparam test_b1_S2043 = 2043;
  localparam test_b1_S2044 = 2044;
  localparam test_b1_S2045 = 2045;
  localparam test_b1_S2046 = 2046;
  localparam test_b1_S2047 = 2047;
  localparam test_b1_S2048 = 2048;
  localparam test_b1_S2049 = 2049;
  localparam test_b1_S2050 = 2050;
  localparam test_b1_S2051 = 2051;
  localparam test_b1_S2052 = 2052;
  localparam test_b1_S2053 = 2053;
  localparam test_b1_S2054 = 2054;
  localparam test_b1_S2055 = 2055;
  localparam test_b1_S2056 = 2056;
  localparam test_b1_S2057 = 2057;
  localparam test_b1_S2058 = 2058;
  localparam test_b1_S2059 = 2059;
  localparam test_b1_S2060 = 2060;
  localparam test_b1_S2061 = 2061;
  localparam test_b1_S2062 = 2062;
  localparam test_b1_S2063 = 2063;
  localparam test_b1_S2064 = 2064;
  localparam test_b1_S2065 = 2065;
  localparam test_b1_S2066 = 2066;
  localparam test_b1_S2067 = 2067;
  localparam test_b1_S2068 = 2068;
  localparam test_b1_S2069 = 2069;
  localparam test_b1_S2070 = 2070;
  localparam test_b1_S2071 = 2071;
  localparam test_b1_S2072 = 2072;
  localparam test_b1_S2073 = 2073;
  localparam test_b1_S2074 = 2074;
  localparam test_b1_S2075 = 2075;
  localparam test_b1_S2076 = 2076;
  localparam test_b1_S2077 = 2077;
  localparam test_b1_S2078 = 2078;
  localparam test_b1_S2079 = 2079;
  localparam test_b1_S2080 = 2080;
  localparam test_b1_S2081 = 2081;
  localparam test_b1_S2082 = 2082;
  localparam test_b1_S2083 = 2083;
  localparam test_b1_S2084 = 2084;
  localparam test_b1_S2085 = 2085;
  localparam test_b1_S2086 = 2086;
  localparam test_b1_S2087 = 2087;
  localparam test_b1_S2088 = 2088;
  localparam test_b1_S2089 = 2089;
  localparam test_b1_S2090 = 2090;
  localparam test_b1_S2091 = 2091;
  localparam test_b1_S2092 = 2092;
  localparam test_b1_S2093 = 2093;
  localparam test_b1_S2094 = 2094;
  localparam test_b1_S2095 = 2095;
  localparam test_b1_S2096 = 2096;
  localparam test_b1_S2097 = 2097;
  localparam test_b1_S2098 = 2098;
  localparam test_b1_S2099 = 2099;
  localparam test_b1_S2100 = 2100;
  localparam test_b1_S2101 = 2101;
  localparam test_b1_S2102 = 2102;
  localparam test_b1_S2103 = 2103;
  localparam test_b1_S2104 = 2104;
  localparam test_b1_S2105 = 2105;
  localparam test_b1_S2106 = 2106;
  localparam test_b1_S2107 = 2107;
  localparam test_b1_S2108 = 2108;
  localparam test_b1_S2109 = 2109;
  localparam test_b1_S2110 = 2110;
  localparam test_b1_S2111 = 2111;
  localparam test_b1_S2112 = 2112;
  localparam test_b1_S2113 = 2113;
  localparam test_b1_S2114 = 2114;
  localparam test_b1_S2115 = 2115;
  localparam test_b1_S2116 = 2116;
  localparam test_b1_S2117 = 2117;
  localparam test_b1_S2118 = 2118;
  localparam test_b1_S2119 = 2119;
  localparam test_b1_S2120 = 2120;
  localparam test_b1_S2121 = 2121;
  localparam test_b1_S2122 = 2122;
  localparam test_b1_S2123 = 2123;
  localparam test_b1_S2124 = 2124;
  localparam test_b1_S2125 = 2125;
  localparam test_b1_S2126 = 2126;
  localparam test_b1_S2127 = 2127;
  localparam test_b1_S2128 = 2128;
  localparam test_b1_S2129 = 2129;
  localparam test_b1_S2130 = 2130;
  localparam test_b1_S2131 = 2131;
  localparam test_b1_S2132 = 2132;
  localparam test_b1_S2133 = 2133;
  localparam test_b1_S2134 = 2134;
  localparam test_b1_S2135 = 2135;
  localparam test_b1_S2136 = 2136;
  localparam test_b1_S2137 = 2137;
  localparam test_b1_S2138 = 2138;
  localparam test_b1_S2139 = 2139;
  localparam test_b1_S2140 = 2140;
  localparam test_b1_S2141 = 2141;
  localparam test_b1_S2142 = 2142;
  localparam test_b1_S2143 = 2143;
  localparam test_b1_S2144 = 2144;
  localparam test_b1_S2145 = 2145;
  localparam test_b1_S2146 = 2146;
  localparam test_b1_S2147 = 2147;
  localparam test_b1_S2148 = 2148;
  localparam test_b1_S2149 = 2149;
  localparam test_b1_S2150 = 2150;
  localparam test_b1_S2151 = 2151;
  localparam test_b1_S2152 = 2152;
  localparam test_b1_S2153 = 2153;
  localparam test_b1_S2154 = 2154;
  localparam test_b1_S2155 = 2155;
  localparam test_b1_S2156 = 2156;
  localparam test_b1_S2157 = 2157;
  localparam test_b1_S2158 = 2158;
  localparam test_b1_S2159 = 2159;
  localparam test_b1_S2160 = 2160;
  localparam test_b1_S2161 = 2161;
  localparam test_b1_S2162 = 2162;
  localparam test_b1_S2163 = 2163;
  localparam test_b1_S2164 = 2164;
  localparam test_b1_S2165 = 2165;
  localparam test_b1_S2166 = 2166;
  localparam test_b1_S2167 = 2167;
  localparam test_b1_S2168 = 2168;
  localparam test_b1_S2169 = 2169;
  localparam test_b1_S2170 = 2170;
  localparam test_b1_S2171 = 2171;
  localparam test_b1_S2172 = 2172;
  localparam test_b1_S2173 = 2173;
  localparam test_b1_S2174 = 2174;
  localparam test_b1_S2175 = 2175;
  localparam test_b1_S2176 = 2176;
  localparam test_b1_S2177 = 2177;
  localparam test_b1_S2178 = 2178;
  localparam test_b1_S2179 = 2179;
  localparam test_b1_S2180 = 2180;
  localparam test_b1_S2181 = 2181;
  localparam test_b1_S2182 = 2182;
  localparam test_b1_S2183 = 2183;
  localparam test_b1_S2184 = 2184;
  localparam test_b1_S2185 = 2185;
  localparam test_b1_S2186 = 2186;
  localparam test_b1_S2187 = 2187;
  localparam test_b1_S2188 = 2188;
  localparam test_b1_S2189 = 2189;
  localparam test_b1_S2190 = 2190;
  localparam test_b1_S2191 = 2191;
  localparam test_b1_S2192 = 2192;
  localparam test_b1_S2193 = 2193;
  localparam test_b1_S2194 = 2194;
  localparam test_b1_S2195 = 2195;
  localparam test_b1_S2196 = 2196;
  localparam test_b1_S2197 = 2197;
  localparam test_b1_S2198 = 2198;
  localparam test_b1_S2199 = 2199;
  localparam test_b1_S2200 = 2200;
  localparam test_b1_S2201 = 2201;
  localparam test_b1_S2202 = 2202;
  localparam test_b1_S2203 = 2203;
  localparam test_b1_S2204 = 2204;
  localparam test_b1_S2205 = 2205;
  localparam test_b1_S2206 = 2206;
  localparam test_b1_S2207 = 2207;
  localparam test_b1_S2208 = 2208;
  localparam test_b1_S2209 = 2209;
  localparam test_b1_S2210 = 2210;
  localparam test_b1_S2211 = 2211;
  localparam test_b1_S2212 = 2212;
  localparam test_b1_S2213 = 2213;
  localparam test_b1_S2214 = 2214;
  localparam test_b1_S2215 = 2215;
  localparam test_b1_S2216 = 2216;
  localparam test_b1_S2217 = 2217;
  localparam test_b1_S2218 = 2218;
  localparam test_b1_S2219 = 2219;
  localparam test_b1_S2220 = 2220;
  localparam test_b1_S2221 = 2221;
  localparam test_b1_S2222 = 2222;
  localparam test_b1_S2223 = 2223;
  localparam test_b1_S2224 = 2224;
  localparam test_b1_S2225 = 2225;
  localparam test_b1_S2226 = 2226;
  localparam test_b1_S2227 = 2227;
  localparam test_b1_S2228 = 2228;
  localparam test_b1_S2229 = 2229;
  localparam test_b1_S2230 = 2230;
  localparam test_b1_S2231 = 2231;
  localparam test_b1_S2232 = 2232;
  localparam test_b1_S2233 = 2233;
  localparam test_b1_S2234 = 2234;
  localparam test_b1_S2235 = 2235;
  localparam test_b1_S2236 = 2236;
  localparam test_b1_S2237 = 2237;
  localparam test_b1_S2238 = 2238;
  localparam test_b1_S2239 = 2239;
  localparam test_b1_S2240 = 2240;
  localparam test_b1_S2241 = 2241;
  localparam test_b1_S2242 = 2242;
  localparam test_b1_S2243 = 2243;
  localparam test_b1_S2244 = 2244;
  localparam test_b1_S2245 = 2245;
  localparam test_b1_S2246 = 2246;
  localparam test_b1_S2247 = 2247;
  localparam test_b1_S2248 = 2248;
  localparam test_b1_S2249 = 2249;
  localparam test_b1_S2250 = 2250;
  localparam test_b1_S2251 = 2251;
  localparam test_b1_S2252 = 2252;
  localparam test_b1_S2253 = 2253;
  localparam test_b1_S2254 = 2254;
  localparam test_b1_S2255 = 2255;
  localparam test_b1_S2256 = 2256;
  localparam test_b1_S2257 = 2257;
  localparam test_b1_S2258 = 2258;
  localparam test_b1_S2259 = 2259;
  localparam test_b1_S2260 = 2260;
  localparam test_b1_S2261 = 2261;
  localparam test_b1_S2262 = 2262;
  localparam test_b1_S2263 = 2263;
  localparam test_b1_S2264 = 2264;
  localparam test_b1_S2265 = 2265;
  localparam test_b1_S2266 = 2266;
  localparam test_b1_S2267 = 2267;
  localparam test_b1_S2268 = 2268;
  localparam test_b1_S2269 = 2269;
  localparam test_b1_S2270 = 2270;
  localparam test_b1_S2271 = 2271;
  localparam test_b1_S2272 = 2272;
  localparam test_b1_S2273 = 2273;
  localparam test_b1_S2274 = 2274;
  localparam test_b1_S2275 = 2275;
  localparam test_b1_S2276 = 2276;
  localparam test_b1_S2277 = 2277;
  localparam test_b1_S2278 = 2278;
  localparam test_b1_S2279 = 2279;
  localparam test_b1_S2280 = 2280;
  localparam test_b1_S2281 = 2281;
  localparam test_b1_S2282 = 2282;
  localparam test_b1_S2283 = 2283;
  localparam test_b1_S2284 = 2284;
  localparam test_b1_S2285 = 2285;
  localparam test_b1_S2286 = 2286;
  localparam test_b1_S2287 = 2287;
  localparam test_b1_S2288 = 2288;
  localparam test_b1_S2289 = 2289;
  localparam test_b1_S2290 = 2290;
  localparam test_b1_S2291 = 2291;
  localparam test_b1_S2292 = 2292;
  localparam test_b1_S2293 = 2293;
  localparam test_b1_S2294 = 2294;
  localparam test_b1_S2295 = 2295;
  localparam test_b1_S2296 = 2296;
  localparam test_b1_S2297 = 2297;
  localparam test_b1_S2298 = 2298;
  localparam test_b1_S2299 = 2299;
  localparam test_b1_S2300 = 2300;
  localparam test_b1_S2301 = 2301;
  localparam test_b1_S2302 = 2302;
  localparam test_b1_S2303 = 2303;
  localparam test_b1_S2304 = 2304;
  localparam test_b1_S2305 = 2305;
  localparam test_b1_S2306 = 2306;
  localparam test_b1_S2307 = 2307;
  localparam test_b1_S2308 = 2308;
  localparam test_b1_S2309 = 2309;
  localparam test_b1_S2310 = 2310;
  localparam test_b1_S2311 = 2311;
  localparam test_b1_S2312 = 2312;
  localparam test_b1_S2313 = 2313;
  localparam test_b1_S2314 = 2314;
  localparam test_b1_S2315 = 2315;
  localparam test_b1_S2316 = 2316;
  localparam test_b1_S2317 = 2317;
  localparam test_b1_S2318 = 2318;
  localparam test_b1_S2319 = 2319;
  localparam test_b1_S2320 = 2320;
  localparam test_b1_S2321 = 2321;
  localparam test_b1_S2322 = 2322;
  localparam test_b1_S2323 = 2323;
  localparam test_b1_S2324 = 2324;
  localparam test_b1_S2325 = 2325;
  localparam test_b1_S2326 = 2326;
  localparam test_b1_S2327 = 2327;
  localparam test_b1_S2328 = 2328;
  localparam test_b1_S2329 = 2329;
  localparam test_b1_S2330 = 2330;
  localparam test_b1_S2331 = 2331;
  localparam test_b1_S2332 = 2332;
  localparam test_b1_S2333 = 2333;
  localparam test_b1_S2334 = 2334;
  localparam test_b1_S2335 = 2335;
  localparam test_b1_S2336 = 2336;
  localparam test_b1_S2337 = 2337;
  localparam test_b1_S2338 = 2338;
  localparam test_b1_S2339 = 2339;
  localparam test_b1_S2340 = 2340;
  localparam test_b1_S2341 = 2341;
  localparam test_b1_S2342 = 2342;
  localparam test_b1_S2343 = 2343;
  localparam test_b1_S2344 = 2344;
  localparam test_b1_S2345 = 2345;
  localparam test_b1_S2346 = 2346;
  localparam test_b1_S2347 = 2347;
  localparam test_b1_S2348 = 2348;
  localparam test_b1_S2349 = 2349;
  localparam test_b1_S2350 = 2350;
  localparam test_b1_S2351 = 2351;
  localparam test_b1_S2352 = 2352;
  localparam test_b1_S2353 = 2353;
  localparam test_b1_S2354 = 2354;
  localparam test_b1_S2355 = 2355;
  localparam test_b1_S2356 = 2356;
  localparam test_b1_S2357 = 2357;
  localparam test_b1_S2358 = 2358;
  localparam test_b1_S2359 = 2359;
  localparam test_b1_S2360 = 2360;
  localparam test_b1_S2361 = 2361;
  localparam test_b1_S2362 = 2362;
  localparam test_b1_S2363 = 2363;
  localparam test_b1_S2364 = 2364;
  localparam test_b1_S2365 = 2365;
  localparam test_b1_S2366 = 2366;
  localparam test_b1_S2367 = 2367;
  localparam test_b1_S2368 = 2368;
  localparam test_b1_S2369 = 2369;
  localparam test_b1_S2370 = 2370;
  localparam test_b1_S2371 = 2371;
  localparam test_b1_S2372 = 2372;
  localparam test_b1_S2373 = 2373;
  localparam test_b1_S2374 = 2374;
  localparam test_b1_S2375 = 2375;
  localparam test_b1_S2376 = 2376;
  localparam test_b1_S2377 = 2377;
  localparam test_b1_S2378 = 2378;
  localparam test_b1_S2379 = 2379;
  localparam test_b1_S2380 = 2380;
  localparam test_b1_S2381 = 2381;
  localparam test_b1_S2382 = 2382;
  localparam test_b1_S2383 = 2383;
  localparam test_b1_S2384 = 2384;
  localparam test_b1_S2385 = 2385;
  localparam test_b1_S2386 = 2386;
  localparam test_b1_S2387 = 2387;
  localparam test_b1_S2388 = 2388;
  localparam test_b1_S2389 = 2389;
  localparam test_b1_S2390 = 2390;
  localparam test_b1_S2391 = 2391;
  localparam test_b1_S2392 = 2392;
  localparam test_b1_S2393 = 2393;
  localparam test_b1_S2394 = 2394;
  localparam test_b1_S2395 = 2395;
  localparam test_b1_S2396 = 2396;
  localparam test_b1_S2397 = 2397;
  localparam test_b1_S2398 = 2398;
  localparam test_b1_S2399 = 2399;
  localparam test_b1_S2400 = 2400;
  localparam test_b1_S2401 = 2401;
  localparam test_b1_S2402 = 2402;
  localparam test_b1_S2403 = 2403;
  localparam test_b1_S2404 = 2404;
  localparam test_b1_S2405 = 2405;
  localparam test_b1_S2406 = 2406;
  localparam test_b1_S2407 = 2407;
  localparam test_b1_S2408 = 2408;
  localparam test_b1_S2409 = 2409;
  localparam test_b1_S2410 = 2410;
  localparam test_b1_S2411 = 2411;
  localparam test_b1_S2412 = 2412;
  localparam test_b1_S2413 = 2413;
  localparam test_b1_S2414 = 2414;
  localparam test_b1_S2415 = 2415;
  localparam test_b1_S2416 = 2416;
  localparam test_b1_S2417 = 2417;
  localparam test_b1_S2418 = 2418;
  localparam test_b1_S2419 = 2419;
  localparam test_b1_S2420 = 2420;
  localparam test_b1_S2421 = 2421;
  localparam test_b1_S2422 = 2422;
  localparam test_b1_S2423 = 2423;
  localparam test_b1_S2424 = 2424;
  localparam test_b1_S2425 = 2425;
  localparam test_b1_S2426 = 2426;
  localparam test_b1_S2427 = 2427;
  localparam test_b1_S2428 = 2428;
  localparam test_b1_S2429 = 2429;
  localparam test_b1_S2430 = 2430;
  localparam test_b1_S2431 = 2431;
  localparam test_b1_S2432 = 2432;
  localparam test_b1_S2433 = 2433;
  localparam test_b1_S2434 = 2434;
  localparam test_b1_S2435 = 2435;
  localparam test_b1_S2436 = 2436;
  localparam test_b1_S2437 = 2437;
  localparam test_b1_S2438 = 2438;
  localparam test_b1_S2439 = 2439;
  localparam test_b1_S2440 = 2440;
  localparam test_b1_S2441 = 2441;
  localparam test_b1_S2442 = 2442;
  localparam test_b1_S2443 = 2443;
  localparam test_b1_S2444 = 2444;
  localparam test_b1_S2445 = 2445;
  localparam test_b1_S2446 = 2446;
  localparam test_b1_S2447 = 2447;
  localparam test_b1_S2448 = 2448;
  localparam test_b1_S2449 = 2449;
  localparam test_b1_S2450 = 2450;
  localparam test_b1_S2451 = 2451;
  localparam test_b1_S2452 = 2452;
  localparam test_b1_S2453 = 2453;
  localparam test_b1_S2454 = 2454;
  localparam test_b1_S2455 = 2455;
  localparam test_b1_S2456 = 2456;
  localparam test_b1_S2457 = 2457;
  localparam test_b1_S2458 = 2458;
  localparam test_b1_S2459 = 2459;
  localparam test_b1_S2460 = 2460;
  localparam test_b1_S2461 = 2461;
  localparam test_b1_S2462 = 2462;
  localparam test_b1_S2463 = 2463;
  localparam test_b1_S2464 = 2464;
  localparam test_b1_S2465 = 2465;
  localparam test_b1_S2466 = 2466;
  localparam test_b1_S2467 = 2467;
  localparam test_b1_S2468 = 2468;
  localparam test_b1_S2469 = 2469;
  localparam test_b1_S2470 = 2470;
  localparam test_b1_S2471 = 2471;
  localparam test_b1_S2472 = 2472;
  localparam test_b1_S2473 = 2473;
  localparam test_b1_S2474 = 2474;
  localparam test_b1_S2475 = 2475;
  localparam test_b1_S2476 = 2476;
  localparam test_b1_S2477 = 2477;
  localparam test_b1_S2478 = 2478;
  localparam test_b1_S2479 = 2479;
  localparam test_b1_S2480 = 2480;
  localparam test_b1_S2481 = 2481;
  localparam test_b1_S2482 = 2482;
  localparam test_b1_S2483 = 2483;
  localparam test_b1_S2484 = 2484;
  localparam test_b1_S2485 = 2485;
  localparam test_b1_S2486 = 2486;
  localparam test_b1_S2487 = 2487;
  localparam test_b1_S2488 = 2488;
  localparam test_b1_S2489 = 2489;
  localparam test_b1_S2490 = 2490;
  localparam test_b1_S2491 = 2491;
  localparam test_b1_S2492 = 2492;
  localparam test_b1_S2493 = 2493;
  localparam test_b1_S2494 = 2494;
  localparam test_b1_S2495 = 2495;
  localparam test_b1_S2496 = 2496;
  localparam test_b1_S2497 = 2497;
  localparam test_b1_S2498 = 2498;
  localparam test_b1_S2499 = 2499;
  localparam test_b1_S2500 = 2500;
  localparam test_b1_S2501 = 2501;
  localparam test_b1_S2502 = 2502;
  localparam test_b1_S2503 = 2503;
  localparam test_b1_S2504 = 2504;
  localparam test_b1_S2505 = 2505;
  localparam test_b1_S2506 = 2506;
  localparam test_b1_S2507 = 2507;
  localparam test_b1_S2508 = 2508;
  localparam test_b1_S2509 = 2509;
  localparam test_b1_S2510 = 2510;
  localparam test_b1_S2511 = 2511;
  localparam test_b1_S2512 = 2512;
  localparam test_b1_S2513 = 2513;
  localparam test_b1_S2514 = 2514;
  localparam test_b1_S2515 = 2515;
  localparam test_b1_S2516 = 2516;
  localparam test_b1_S2517 = 2517;
  localparam test_b1_S2518 = 2518;
  localparam test_b1_S2519 = 2519;
  localparam test_b1_S2520 = 2520;
  localparam test_b1_S2521 = 2521;
  localparam test_b1_S2522 = 2522;
  localparam test_b1_S2523 = 2523;
  localparam test_b1_S2524 = 2524;
  localparam test_b1_S2525 = 2525;
  localparam test_b1_S2526 = 2526;
  localparam test_b1_S2527 = 2527;
  localparam test_b1_S2528 = 2528;
  localparam test_b1_S2529 = 2529;
  localparam test_b1_S2530 = 2530;
  localparam test_b1_S2531 = 2531;
  localparam test_b1_S2532 = 2532;
  localparam test_b1_S2533 = 2533;
  localparam test_b1_S2534 = 2534;
  localparam test_b1_S2535 = 2535;
  localparam test_b1_S2536 = 2536;
  localparam test_b1_S2537 = 2537;
  localparam test_b1_S2538 = 2538;
  localparam test_b1_S2539 = 2539;
  localparam test_b1_S2540 = 2540;
  localparam test_b1_S2541 = 2541;
  localparam test_b1_S2542 = 2542;
  localparam test_b1_S2543 = 2543;
  localparam test_b1_S2544 = 2544;
  localparam test_b1_S2545 = 2545;
  localparam test_b1_S2546 = 2546;
  localparam test_b1_S2547 = 2547;
  localparam test_b1_S2548 = 2548;
  localparam test_b1_S2549 = 2549;
  localparam test_b1_S2550 = 2550;
  localparam test_b1_S2551 = 2551;
  localparam test_b1_S2552 = 2552;
  localparam test_b1_S2553 = 2553;
  localparam test_b1_S2554 = 2554;
  localparam test_b1_S2555 = 2555;
  localparam test_b1_S2556 = 2556;
  localparam test_b1_S2557 = 2557;
  localparam test_b1_S2558 = 2558;
  localparam test_b1_S2559 = 2559;
  localparam test_b1_S2560 = 2560;
  localparam test_b1_S2561 = 2561;
  localparam test_b1_S2562 = 2562;
  localparam test_b1_S2563 = 2563;
  localparam test_b1_S2564 = 2564;
  localparam test_b1_S2565 = 2565;
  localparam test_b1_S2566 = 2566;
  localparam test_b1_S2567 = 2567;
  localparam test_b1_S2568 = 2568;
  localparam test_b1_S2569 = 2569;
  localparam test_b1_S2570 = 2570;
  localparam test_b1_S2571 = 2571;
  localparam test_b1_S2572 = 2572;
  localparam test_b1_S2573 = 2573;
  localparam test_b1_S2574 = 2574;
  localparam test_b1_S2575 = 2575;
  localparam test_b1_S2576 = 2576;
  localparam test_b1_S2577 = 2577;
  localparam test_b1_S2578 = 2578;
  localparam test_b1_S2579 = 2579;
  localparam test_b1_S2580 = 2580;
  localparam test_b1_S2581 = 2581;
  localparam test_b1_S2582 = 2582;
  localparam test_b1_S2583 = 2583;
  localparam test_b1_S2584 = 2584;
  localparam test_b1_S2585 = 2585;
  localparam test_b1_S2586 = 2586;
  localparam test_b1_S2587 = 2587;
  localparam test_b1_S2588 = 2588;
  localparam test_b1_S2589 = 2589;
  localparam test_b1_S2590 = 2590;
  localparam test_b1_S2591 = 2591;
  localparam test_b1_S2592 = 2592;
  localparam test_b1_S2593 = 2593;
  localparam test_b1_S2594 = 2594;
  localparam test_b1_S2595 = 2595;
  localparam test_b1_S2596 = 2596;
  localparam test_b1_S2597 = 2597;
  localparam test_b1_S2598 = 2598;
  localparam test_b1_S2599 = 2599;
  localparam test_b1_S2600 = 2600;
  localparam test_b1_S2601 = 2601;
  localparam test_b1_S2602 = 2602;
  localparam test_b1_S2603 = 2603;
  localparam test_b1_S2604 = 2604;
  localparam test_b1_S2605 = 2605;
  localparam test_b1_S2606 = 2606;
  localparam test_b1_S2607 = 2607;
  localparam test_b1_S2608 = 2608;
  localparam test_b1_S2609 = 2609;
  localparam test_b1_S2610 = 2610;
  localparam test_b1_S2611 = 2611;
  localparam test_b1_S2612 = 2612;
  localparam test_b1_S2613 = 2613;
  localparam test_b1_S2614 = 2614;
  localparam test_b1_S2615 = 2615;
  localparam test_b1_S2616 = 2616;
  localparam test_b1_S2617 = 2617;
  localparam test_b1_S2618 = 2618;
  localparam test_b1_S2619 = 2619;
  localparam test_b1_S2620 = 2620;
  localparam test_b1_S2621 = 2621;
  localparam test_b1_S2622 = 2622;
  localparam test_b1_S2623 = 2623;
  localparam test_b1_S2624 = 2624;
  localparam test_b1_S2625 = 2625;
  localparam test_b1_S2626 = 2626;
  localparam test_b1_S2627 = 2627;
  localparam test_b1_S2628 = 2628;
  localparam test_b1_S2629 = 2629;
  localparam test_b1_S2630 = 2630;
  localparam test_b1_S2631 = 2631;
  localparam test_b1_S2632 = 2632;
  localparam test_b1_S2633 = 2633;
  localparam test_b1_S2634 = 2634;
  localparam test_b1_S2635 = 2635;
  localparam test_b1_S2636 = 2636;
  localparam test_b1_S2637 = 2637;
  localparam test_b1_S2638 = 2638;
  localparam test_b1_S2639 = 2639;
  localparam test_b1_S2640 = 2640;
  localparam test_b1_S2641 = 2641;
  localparam test_b1_S2642 = 2642;
  localparam test_b1_S2643 = 2643;
  localparam test_b1_S2644 = 2644;
  localparam test_b1_S2645 = 2645;
  localparam test_b1_S2646 = 2646;
  localparam test_b1_S2647 = 2647;
  localparam test_b1_S2648 = 2648;
  localparam test_b1_S2649 = 2649;
  localparam test_b1_S2650 = 2650;
  localparam test_b1_S2651 = 2651;
  localparam test_b1_S2652 = 2652;
  localparam test_b1_S2653 = 2653;
  localparam test_b1_S2654 = 2654;
  localparam test_b1_S2655 = 2655;
  localparam test_b1_S2656 = 2656;
  localparam test_b1_S2657 = 2657;
  localparam test_b1_S2658 = 2658;
  localparam test_b1_S2659 = 2659;
  localparam test_b1_S2660 = 2660;
  localparam test_b1_S2661 = 2661;
  localparam test_b1_S2662 = 2662;
  localparam test_b1_S2663 = 2663;
  localparam test_b1_S2664 = 2664;
  localparam test_b1_S2665 = 2665;
  localparam test_b1_S2666 = 2666;
  localparam test_b1_S2667 = 2667;
  localparam test_b1_S2668 = 2668;
  localparam test_b1_S2669 = 2669;
  localparam test_b1_S2670 = 2670;
  localparam test_b1_S2671 = 2671;
  localparam test_b1_S2672 = 2672;
  localparam test_b1_S2673 = 2673;
  localparam test_b1_S2674 = 2674;
  localparam test_b1_S2675 = 2675;
  localparam test_b1_S2676 = 2676;
  localparam test_b1_S2677 = 2677;
  localparam test_b1_S2678 = 2678;
  localparam test_b1_S2679 = 2679;
  localparam test_b1_S2680 = 2680;
  localparam test_b1_S2681 = 2681;
  localparam test_b1_S2682 = 2682;
  localparam test_b1_S2683 = 2683;
  localparam test_b1_S2684 = 2684;
  localparam test_b1_S2685 = 2685;
  localparam test_b1_S2686 = 2686;
  localparam test_b1_S2687 = 2687;
  localparam test_b1_S2688 = 2688;
  localparam test_b1_S2689 = 2689;
  localparam test_b1_S2690 = 2690;
  localparam test_b1_S2691 = 2691;
  localparam test_b1_S2692 = 2692;
  localparam test_b1_S2693 = 2693;
  localparam test_b1_S2694 = 2694;
  localparam test_b1_S2695 = 2695;
  localparam test_b1_S2696 = 2696;
  localparam test_b1_S2697 = 2697;
  localparam test_b1_S2698 = 2698;
  localparam test_b1_S2699 = 2699;
  localparam test_b1_S2700 = 2700;
  localparam test_b1_S2701 = 2701;
  localparam test_b1_S2702 = 2702;
  localparam test_b1_S2703 = 2703;
  localparam test_b1_S2704 = 2704;
  localparam test_b1_S2705 = 2705;
  localparam test_b1_S2706 = 2706;
  localparam test_b1_S2707 = 2707;
  localparam test_b1_S2708 = 2708;
  localparam test_b1_S2709 = 2709;
  localparam test_b1_S2710 = 2710;
  localparam test_b1_S2711 = 2711;
  localparam test_b1_S2712 = 2712;
  localparam test_b1_S2713 = 2713;
  localparam test_b1_S2714 = 2714;
  localparam test_b1_S2715 = 2715;
  localparam test_b1_S2716 = 2716;
  localparam test_b1_S2717 = 2717;
  localparam test_b1_S2718 = 2718;
  localparam test_b1_S2719 = 2719;
  localparam test_b1_S2720 = 2720;
  localparam test_b1_S2721 = 2721;
  localparam test_b1_S2722 = 2722;
  localparam test_b1_S2723 = 2723;
  localparam test_b1_S2724 = 2724;
  localparam test_b1_S2725 = 2725;
  localparam test_b1_S2726 = 2726;
  localparam test_b1_S2727 = 2727;
  localparam test_b1_S2728 = 2728;
  localparam test_b1_S2729 = 2729;
  localparam test_b1_S2730 = 2730;
  localparam test_b1_S2731 = 2731;
  localparam test_b1_S2732 = 2732;
  localparam test_b1_S2733 = 2733;
  localparam test_b1_S2734 = 2734;
  localparam test_b1_S2735 = 2735;
  localparam test_b1_S2736 = 2736;
  localparam test_b1_S2737 = 2737;
  localparam test_b1_S2738 = 2738;
  localparam test_b1_S2739 = 2739;
  localparam test_b1_S2740 = 2740;
  localparam test_b1_S2741 = 2741;
  localparam test_b1_S2742 = 2742;
  localparam test_b1_S2743 = 2743;
  localparam test_b1_S2744 = 2744;
  localparam test_b1_S2745 = 2745;
  localparam test_b1_S2746 = 2746;
  localparam test_b1_S2747 = 2747;
  localparam test_b1_S2748 = 2748;
  localparam test_b1_S2749 = 2749;
  localparam test_b1_S2750 = 2750;
  localparam test_b1_S2751 = 2751;
  localparam test_b1_S2752 = 2752;
  localparam test_b1_S2753 = 2753;
  localparam test_b1_S2754 = 2754;
  localparam test_b1_S2755 = 2755;
  localparam test_b1_S2756 = 2756;
  localparam test_b1_S2757 = 2757;
  localparam test_b1_S2758 = 2758;
  localparam test_b1_S2759 = 2759;
  localparam test_b1_S2760 = 2760;
  localparam test_b1_S2761 = 2761;
  localparam test_b1_S2762 = 2762;
  localparam test_b1_S2763 = 2763;
  localparam test_b1_S2764 = 2764;
  localparam test_b1_S2765 = 2765;
  localparam test_b1_S2766 = 2766;
  localparam test_b1_S2767 = 2767;
  localparam test_b1_S2768 = 2768;
  localparam test_b1_S2769 = 2769;
  localparam test_b1_S2770 = 2770;
  localparam test_b1_S2771 = 2771;
  localparam test_b1_S2772 = 2772;
  localparam test_b1_S2773 = 2773;
  localparam test_b1_S2774 = 2774;
  localparam test_b1_S2775 = 2775;
  localparam test_b1_S2776 = 2776;
  localparam test_b1_S2777 = 2777;
  localparam test_b1_S2778 = 2778;
  localparam test_b1_S2779 = 2779;
  localparam test_b1_S2780 = 2780;
  localparam test_b1_S2781 = 2781;
  localparam test_b1_S2782 = 2782;
  localparam test_b1_S2783 = 2783;
  localparam test_b1_S2784 = 2784;
  localparam test_b1_S2785 = 2785;
  localparam test_b1_S2786 = 2786;
  localparam test_b1_S2787 = 2787;
  localparam test_b1_S2788 = 2788;
  localparam test_b1_S2789 = 2789;
  localparam test_b1_S2790 = 2790;
  localparam test_b1_S2791 = 2791;
  localparam test_b1_S2792 = 2792;
  localparam test_b1_S2793 = 2793;
  localparam test_b1_S2794 = 2794;
  localparam test_b1_S2795 = 2795;
  localparam test_b1_S2796 = 2796;
  localparam test_b1_S2797 = 2797;
  localparam test_b1_S2798 = 2798;
  localparam test_b1_S2799 = 2799;
  localparam test_b1_S2800 = 2800;
  localparam test_b1_S2801 = 2801;
  localparam test_b1_S2802 = 2802;
  localparam test_b1_S2803 = 2803;
  localparam test_b1_S2804 = 2804;
  localparam test_b1_S2805 = 2805;
  localparam test_b1_S2806 = 2806;
  localparam test_b1_S2807 = 2807;
  localparam test_b1_S2808 = 2808;
  localparam test_b1_S2809 = 2809;
  localparam test_b1_S2810 = 2810;
  localparam test_b1_S2811 = 2811;
  localparam test_b1_S2812 = 2812;
  localparam test_b1_S2813 = 2813;
  localparam test_b1_S2814 = 2814;
  localparam test_b1_S2815 = 2815;
  localparam test_b1_S2816 = 2816;
  localparam test_b1_S2817 = 2817;
  localparam test_b1_S2818 = 2818;
  localparam test_b1_S2819 = 2819;
  localparam test_b1_S2820 = 2820;
  localparam test_b1_S2821 = 2821;
  localparam test_b1_S2822 = 2822;
  localparam test_b1_S2823 = 2823;
  localparam test_b1_S2824 = 2824;
  localparam test_b1_S2825 = 2825;
  localparam test_b1_S2826 = 2826;
  localparam test_b1_S2827 = 2827;
  localparam test_b1_S2828 = 2828;
  localparam test_b1_S2829 = 2829;
  localparam test_b1_S2830 = 2830;
  localparam test_b1_S2831 = 2831;
  localparam test_b1_S2832 = 2832;
  localparam test_b1_S2833 = 2833;
  localparam test_b1_S2834 = 2834;
  localparam test_b1_S2835 = 2835;
  localparam test_b1_S2836 = 2836;
  localparam test_b1_S2837 = 2837;
  localparam test_b1_S2838 = 2838;
  localparam test_b1_S2839 = 2839;
  localparam test_b1_S2840 = 2840;
  localparam test_b1_S2841 = 2841;
  localparam test_b1_S2842 = 2842;
  localparam test_b1_S2843 = 2843;
  localparam test_b1_S2844 = 2844;
  localparam test_b1_S2845 = 2845;
  localparam test_b1_S2846 = 2846;
  localparam test_b1_S2847 = 2847;
  localparam test_b1_S2848 = 2848;
  localparam test_b1_S2849 = 2849;
  localparam test_b1_S2850 = 2850;
  localparam test_b1_S2851 = 2851;
  localparam test_b1_S2852 = 2852;
  localparam test_b1_S2853 = 2853;
  localparam test_b1_S2854 = 2854;
  localparam test_b1_S2855 = 2855;
  localparam test_b1_S2856 = 2856;
  localparam test_b1_S2857 = 2857;
  localparam test_b1_S2858 = 2858;
  localparam test_b1_S2859 = 2859;
  localparam test_b1_S2860 = 2860;
  localparam test_b1_S2861 = 2861;
  localparam test_b1_S2862 = 2862;
  localparam test_b1_S2863 = 2863;
  localparam test_b1_S2864 = 2864;
  localparam test_b1_S2865 = 2865;
  localparam test_b1_S2866 = 2866;
  localparam test_b1_S2867 = 2867;
  localparam test_b1_S2868 = 2868;
  localparam test_b1_S2869 = 2869;
  localparam test_b1_S2870 = 2870;
  localparam test_b1_S2871 = 2871;
  localparam test_b1_S2872 = 2872;
  localparam test_b1_S2873 = 2873;
  localparam test_b1_S2874 = 2874;
  localparam test_b1_S2875 = 2875;
  localparam test_b1_S2876 = 2876;
  localparam test_b1_S2877 = 2877;
  localparam test_b1_S2878 = 2878;
  localparam test_b1_S2879 = 2879;
  localparam test_b1_S2880 = 2880;
  localparam test_b1_S2881 = 2881;
  localparam test_b1_S2882 = 2882;
  localparam test_b1_S2883 = 2883;
  localparam test_b1_S2884 = 2884;
  localparam test_b1_S2885 = 2885;
  localparam test_b1_S2886 = 2886;
  localparam test_b1_S2887 = 2887;
  localparam test_b1_S2888 = 2888;
  localparam test_b1_S2889 = 2889;
  localparam test_b1_S2890 = 2890;
  localparam test_b1_S2891 = 2891;
  localparam test_b1_S2892 = 2892;
  localparam test_b1_S2893 = 2893;
  localparam test_b1_S2894 = 2894;
  localparam test_b1_S2895 = 2895;
  localparam test_b1_S2896 = 2896;
  localparam test_b1_S2897 = 2897;
  localparam test_b1_S2898 = 2898;
  localparam test_b1_S2899 = 2899;
  localparam test_b1_S2900 = 2900;
  localparam test_b1_S2901 = 2901;
  localparam test_b1_S2902 = 2902;
  localparam test_b1_S2903 = 2903;
  localparam test_b1_S2904 = 2904;
  localparam test_b1_S2905 = 2905;
  localparam test_b1_S2906 = 2906;
  localparam test_b1_S2907 = 2907;
  localparam test_b1_S2908 = 2908;
  localparam test_b1_S2909 = 2909;
  localparam test_b1_S2910 = 2910;
  localparam test_b1_S2911 = 2911;
  localparam test_b1_S2912 = 2912;
  localparam test_b1_S2913 = 2913;
  localparam test_b1_S2914 = 2914;
  localparam test_b1_S2915 = 2915;
  localparam test_b1_S2916 = 2916;
  localparam test_b1_S2917 = 2917;
  localparam test_b1_S2918 = 2918;
  localparam test_b1_S2919 = 2919;
  localparam test_b1_S2920 = 2920;
  localparam test_b1_S2921 = 2921;
  localparam test_b1_S2922 = 2922;
  localparam test_b1_S2923 = 2923;
  localparam test_b1_S2924 = 2924;
  localparam test_b1_S2925 = 2925;
  localparam test_b1_S2926 = 2926;
  localparam test_b1_S2927 = 2927;
  localparam test_b1_S2928 = 2928;
  localparam test_b1_S2929 = 2929;
  localparam test_b1_S2930 = 2930;
  localparam test_b1_S2931 = 2931;
  localparam test_b1_S2932 = 2932;
  localparam test_b1_S2933 = 2933;
  localparam test_b1_S2934 = 2934;
  localparam test_b1_S2935 = 2935;
  localparam test_b1_S2936 = 2936;
  localparam test_b1_S2937 = 2937;
  localparam test_b1_S2938 = 2938;
  localparam test_b1_S2939 = 2939;
  localparam test_b1_S2940 = 2940;
  localparam test_b1_S2941 = 2941;
  localparam test_b1_S2942 = 2942;
  localparam test_b1_S2943 = 2943;
  localparam test_b1_S2944 = 2944;
  localparam test_b1_S2945 = 2945;
  localparam test_b1_S2946 = 2946;
  localparam test_b1_S2947 = 2947;
  localparam test_b1_S2948 = 2948;
  localparam test_b1_S2949 = 2949;
  localparam test_b1_S2950 = 2950;
  localparam test_b1_S2951 = 2951;
  localparam test_b1_S2952 = 2952;
  localparam test_b1_S2953 = 2953;
  localparam test_b1_S2954 = 2954;
  localparam test_b1_S2955 = 2955;
  localparam test_b1_S2956 = 2956;
  localparam test_b1_S2957 = 2957;
  localparam test_b1_S2958 = 2958;
  localparam test_b1_S2959 = 2959;
  localparam test_b1_S2960 = 2960;
  localparam test_b1_S2961 = 2961;
  localparam test_b1_S2962 = 2962;
  localparam test_b1_S2963 = 2963;
  localparam test_b1_S2964 = 2964;
  localparam test_b1_S2965 = 2965;
  localparam test_b1_S2966 = 2966;
  localparam test_b1_S2967 = 2967;
  localparam test_b1_S2968 = 2968;
  localparam test_b1_S2969 = 2969;
  localparam test_b1_S2970 = 2970;
  localparam test_b1_S2971 = 2971;
  localparam test_b1_S2972 = 2972;
  localparam test_b1_S2973 = 2973;
  localparam test_b1_S2974 = 2974;
  localparam test_b1_S2975 = 2975;
  localparam test_b1_S2976 = 2976;
  localparam test_b1_S2977 = 2977;
  localparam test_b1_S2978 = 2978;
  localparam test_b1_S2979 = 2979;
  localparam test_b1_S2980 = 2980;
  localparam test_b1_S2981 = 2981;
  localparam test_b1_S2982 = 2982;
  localparam test_b1_S2983 = 2983;
  localparam test_b1_S2984 = 2984;
  localparam test_b1_S2985 = 2985;
  localparam test_b1_S2986 = 2986;
  localparam test_b1_S2987 = 2987;
  localparam test_b1_S2988 = 2988;
  localparam test_b1_S2989 = 2989;
  localparam test_b1_S2990 = 2990;
  localparam test_b1_S2991 = 2991;
  localparam test_b1_S2992 = 2992;
  localparam test_b1_S2993 = 2993;
  localparam test_b1_S2994 = 2994;
  localparam test_b1_S2995 = 2995;
  localparam test_b1_S2996 = 2996;
  localparam test_b1_S2997 = 2997;
  localparam test_b1_S2998 = 2998;
  localparam test_b1_S2999 = 2999;
  localparam test_b1_S3000 = 3000;
  localparam test_b1_S3001 = 3001;
  localparam test_b1_S3002 = 3002;
  localparam test_b1_S3003 = 3003;
  localparam test_b1_S3004 = 3004;
  localparam test_b1_S3005 = 3005;
  localparam test_b1_S3006 = 3006;
  localparam test_b1_S3007 = 3007;
  localparam test_b1_S3008 = 3008;
  localparam test_b1_S3009 = 3009;
  localparam test_b1_S3010 = 3010;
  localparam test_b1_S3011 = 3011;
  localparam test_b1_S3012 = 3012;
  localparam test_b1_S3013 = 3013;
  localparam test_b1_S3014 = 3014;
  localparam test_b1_S3015 = 3015;
  localparam test_b1_S3016 = 3016;
  localparam test_b1_S3017 = 3017;
  localparam test_b1_S3018 = 3018;
  localparam test_b1_S3019 = 3019;
  localparam test_b1_S3020 = 3020;
  localparam test_b1_S3021 = 3021;
  localparam test_b1_S3022 = 3022;
  localparam test_b1_S3023 = 3023;
  localparam test_b1_S3024 = 3024;
  localparam test_b1_S3025 = 3025;
  localparam test_b1_S3026 = 3026;
  localparam test_b1_S3027 = 3027;
  localparam test_b1_S3028 = 3028;
  localparam test_b1_S3029 = 3029;
  localparam test_b1_S3030 = 3030;
  localparam test_b1_S3031 = 3031;
  localparam test_b1_S3032 = 3032;
  localparam test_b1_S3033 = 3033;
  localparam test_b1_S3034 = 3034;
  localparam test_b1_S3035 = 3035;
  localparam test_b1_S3036 = 3036;
  localparam test_b1_S3037 = 3037;
  localparam test_b1_S3038 = 3038;
  localparam test_b1_S3039 = 3039;
  localparam test_b1_S3040 = 3040;
  localparam test_b1_S3041 = 3041;
  localparam test_b1_S3042 = 3042;
  localparam test_b1_S3043 = 3043;
  localparam test_b1_S3044 = 3044;
  localparam test_b1_S3045 = 3045;
  localparam test_b1_S3046 = 3046;
  localparam test_b1_S3047 = 3047;
  localparam test_b1_S3048 = 3048;
  localparam test_b1_S3049 = 3049;
  localparam test_b1_S3050 = 3050;
  localparam test_b1_S3051 = 3051;
  localparam test_b1_S3052 = 3052;
  localparam test_b1_S3053 = 3053;
  localparam test_b1_S3054 = 3054;
  localparam test_b1_S3055 = 3055;
  localparam test_b1_S3056 = 3056;
  localparam test_b1_S3057 = 3057;
  localparam test_b1_S3058 = 3058;
  localparam test_b1_S3059 = 3059;
  localparam test_b1_S3060 = 3060;
  localparam test_b1_S3061 = 3061;
  localparam test_b1_S3062 = 3062;
  localparam test_b1_S3063 = 3063;
  localparam test_b1_S3064 = 3064;
  localparam test_b1_S3065 = 3065;
  localparam test_b1_S3066 = 3066;
  localparam test_b1_S3067 = 3067;
  localparam test_b1_S3068 = 3068;
  localparam test_b1_S3069 = 3069;
  localparam test_b1_S3070 = 3070;
  localparam test_b1_S3071 = 3071;
  localparam test_b1_S3072 = 3072;
  localparam test_b1_S3073 = 3073;
  localparam test_b1_S3074 = 3074;
  localparam test_b1_S3075 = 3075;
  localparam test_b1_S3076 = 3076;
  localparam test_b1_S3077 = 3077;
  localparam test_b1_S3078 = 3078;
  localparam test_b1_S3079 = 3079;
  localparam test_b1_S3080 = 3080;
  localparam test_b1_S3081 = 3081;
  localparam test_b1_S3082 = 3082;
  localparam test_b1_S3083 = 3083;
  localparam test_b1_S3084 = 3084;
  localparam test_b1_S3085 = 3085;
  localparam test_b1_S3086 = 3086;
  localparam test_b1_S3087 = 3087;
  localparam test_b1_S3088 = 3088;
  localparam test_b1_S3089 = 3089;
  localparam test_b1_S3090 = 3090;
  localparam test_b1_S3091 = 3091;
  localparam test_b1_S3092 = 3092;
  localparam test_b1_S3093 = 3093;
  localparam test_b1_S3094 = 3094;
  localparam test_b1_S3095 = 3095;
  localparam test_b1_S3096 = 3096;
  localparam test_b1_S3097 = 3097;
  localparam test_b1_S3098 = 3098;
  localparam test_b1_S3099 = 3099;
  localparam test_b1_S3100 = 3100;
  localparam test_b1_S3101 = 3101;
  localparam test_b1_S3102 = 3102;
  localparam test_b1_S3103 = 3103;
  localparam test_b1_S3104 = 3104;
  localparam test_b1_S3105 = 3105;
  localparam test_b1_S3106 = 3106;
  localparam test_b1_S3107 = 3107;
  localparam test_b1_S3108 = 3108;
  localparam test_b1_S3109 = 3109;
  localparam test_b1_S3110 = 3110;
  localparam test_b1_S3111 = 3111;
  localparam test_b1_S3112 = 3112;
  localparam test_b1_S3113 = 3113;
  localparam test_b1_S3114 = 3114;
  localparam test_b1_S3115 = 3115;
  localparam test_b1_S3116 = 3116;
  localparam test_b1_S3117 = 3117;
  localparam test_b1_S3118 = 3118;
  localparam test_b1_S3119 = 3119;
  localparam test_b1_S3120 = 3120;
  localparam test_b1_S3121 = 3121;
  localparam test_b1_S3122 = 3122;
  localparam test_b1_S3123 = 3123;
  localparam test_b1_S3124 = 3124;
  localparam test_b1_S3125 = 3125;
  localparam test_b1_S3126 = 3126;
  localparam test_b1_S3127 = 3127;
  localparam test_b1_S3128 = 3128;
  localparam test_b1_S3129 = 3129;
  localparam test_b1_S3130 = 3130;
  localparam test_b1_S3131 = 3131;
  localparam test_b1_S3132 = 3132;
  localparam test_b1_S3133 = 3133;
  localparam test_b1_S3134 = 3134;
  localparam test_b1_S3135 = 3135;
  localparam test_b1_S3136 = 3136;
  localparam test_b1_S3137 = 3137;
  localparam test_b1_S3138 = 3138;
  localparam test_b1_S3139 = 3139;
  localparam test_b1_S3140 = 3140;
  localparam test_b1_S3141 = 3141;
  localparam test_b1_S3142 = 3142;
  localparam test_b1_S3143 = 3143;
  localparam test_b1_S3144 = 3144;
  localparam test_b1_S3145 = 3145;
  localparam test_b1_S3146 = 3146;
  localparam test_b1_S3147 = 3147;
  localparam test_b1_S3148 = 3148;
  localparam test_b1_S3149 = 3149;
  localparam test_b1_S3150 = 3150;
  localparam test_b1_S3151 = 3151;
  localparam test_b1_S3152 = 3152;
  localparam test_b1_S3153 = 3153;
  localparam test_b1_S3154 = 3154;
  localparam test_b1_S3155 = 3155;
  localparam test_b1_S3156 = 3156;
  localparam test_b1_S3157 = 3157;
  localparam test_b1_S3158 = 3158;
  localparam test_b1_S3159 = 3159;
  localparam test_b1_S3160 = 3160;
  localparam test_b1_S3161 = 3161;
  localparam test_b1_S3162 = 3162;
  localparam test_b1_S3163 = 3163;
  localparam test_b1_S3164 = 3164;
  localparam test_b1_S3165 = 3165;
  localparam test_b1_S3166 = 3166;
  localparam test_b1_S3167 = 3167;
  localparam test_b1_S3168 = 3168;
  localparam test_b1_S3169 = 3169;
  localparam test_b1_S3170 = 3170;
  localparam test_b1_S3171 = 3171;
  localparam test_b1_S3172 = 3172;
  localparam test_b1_S3173 = 3173;
  localparam test_b1_S3174 = 3174;
  localparam test_b1_S3175 = 3175;
  localparam test_b1_S3176 = 3176;
  localparam test_b1_S3177 = 3177;
  localparam test_b1_S3178 = 3178;
  localparam test_b1_S3179 = 3179;
  localparam test_b1_S3180 = 3180;
  localparam test_b1_S3181 = 3181;
  localparam test_b1_S3182 = 3182;
  localparam test_b1_S3183 = 3183;
  localparam test_b1_S3184 = 3184;
  localparam test_b1_S3185 = 3185;
  localparam test_b1_S3186 = 3186;
  localparam test_b1_S3187 = 3187;
  localparam test_b1_S3188 = 3188;
  localparam test_b1_S3189 = 3189;
  localparam test_b1_S3190 = 3190;
  localparam test_b1_S3191 = 3191;
  localparam test_b1_S3192 = 3192;
  localparam test_b1_S3193 = 3193;
  localparam test_b1_S3194 = 3194;
  localparam test_b1_S3195 = 3195;
  localparam test_b1_S3196 = 3196;
  localparam test_b1_S3197 = 3197;
  localparam test_b1_S3198 = 3198;
  localparam test_b1_S3199 = 3199;
  localparam test_b1_S3200 = 3200;
  localparam test_b1_S3201 = 3201;
  localparam test_b1_S3202 = 3202;
  localparam test_b1_S3203 = 3203;
  localparam test_b1_S3204 = 3204;
  localparam test_b1_S3205 = 3205;
  localparam test_b1_S3206 = 3206;
  localparam test_b1_S3207 = 3207;
  localparam test_b1_S3208 = 3208;
  localparam test_b1_S3209 = 3209;
  localparam test_b1_S3210 = 3210;
  localparam test_b1_S3211 = 3211;
  localparam test_b1_S3212 = 3212;
  localparam test_b1_S3213 = 3213;
  localparam test_b1_S3214 = 3214;
  localparam test_b1_S3215 = 3215;
  localparam test_b1_S3216 = 3216;
  localparam test_b1_S3217 = 3217;
  localparam test_b1_S3218 = 3218;
  localparam test_b1_S3219 = 3219;
  localparam test_b1_S3220 = 3220;
  localparam test_b1_S3221 = 3221;
  localparam test_b1_S3222 = 3222;
  localparam test_b1_S3223 = 3223;
  localparam test_b1_S3224 = 3224;
  localparam test_b1_S3225 = 3225;
  localparam test_b1_S3226 = 3226;
  localparam test_b1_S3227 = 3227;
  localparam test_b1_S3228 = 3228;
  localparam test_b1_S3229 = 3229;
  localparam test_b1_S3230 = 3230;
  localparam test_b1_S3231 = 3231;
  localparam test_b1_S3232 = 3232;
  localparam test_b1_S3233 = 3233;
  localparam test_b1_S3234 = 3234;
  localparam test_b1_S3235 = 3235;
  localparam test_b1_S3236 = 3236;
  localparam test_b1_S3237 = 3237;
  localparam test_b1_S3238 = 3238;
  localparam test_b1_S3239 = 3239;
  localparam test_b1_S3240 = 3240;
  localparam test_b1_S3241 = 3241;
  localparam test_b1_S3242 = 3242;
  localparam test_b1_S3243 = 3243;
  localparam test_b1_S3244 = 3244;
  localparam test_b1_S3245 = 3245;
  localparam test_b1_S3246 = 3246;
  localparam test_b1_S3247 = 3247;
  localparam test_b1_S3248 = 3248;
  localparam test_b1_S3249 = 3249;
  localparam test_b1_S3250 = 3250;
  localparam test_b1_S3251 = 3251;
  localparam test_b1_S3252 = 3252;
  localparam test_b1_S3253 = 3253;
  localparam test_b1_S3254 = 3254;
  localparam test_b1_S3255 = 3255;
  localparam test_b1_S3256 = 3256;
  localparam test_b1_S3257 = 3257;
  localparam test_b1_S3258 = 3258;
  localparam test_b1_S3259 = 3259;
  localparam test_b1_S3260 = 3260;
  localparam test_b1_S3261 = 3261;
  localparam test_b1_S3262 = 3262;
  localparam test_b1_S3263 = 3263;
  localparam test_b1_S3264 = 3264;
  localparam test_b1_S3265 = 3265;
  localparam test_b1_S3266 = 3266;
  localparam test_b1_S3267 = 3267;
  localparam test_b1_S3268 = 3268;
  localparam test_b1_S3269 = 3269;
  localparam test_b1_S3270 = 3270;
  localparam test_b1_S3271 = 3271;
  localparam test_b1_S3272 = 3272;
  localparam test_b1_S3273 = 3273;
  localparam test_b1_S3274 = 3274;
  localparam test_b1_S3275 = 3275;
  localparam test_b1_S3276 = 3276;
  localparam test_b1_S3277 = 3277;
  localparam test_b1_S3278 = 3278;
  localparam test_b1_S3279 = 3279;
  localparam test_b1_S3280 = 3280;
  localparam test_b1_S3281 = 3281;
  localparam test_b1_S3282 = 3282;
  localparam test_b1_S3283 = 3283;
  localparam test_b1_S3284 = 3284;
  localparam test_b1_S3285 = 3285;
  localparam test_b1_S3286 = 3286;
  localparam test_b1_S3287 = 3287;
  localparam test_b1_S3288 = 3288;
  localparam test_b1_S3289 = 3289;
  localparam test_b1_S3290 = 3290;
  localparam test_b1_S3291 = 3291;
  localparam test_b1_S3292 = 3292;
  localparam test_b1_S3293 = 3293;
  localparam test_b1_S3294 = 3294;
  localparam test_b1_S3295 = 3295;
  localparam test_b1_S3296 = 3296;
  localparam test_b1_S3297 = 3297;
  localparam test_b1_S3298 = 3298;
  localparam test_b1_S3299 = 3299;
  localparam test_b1_S3300 = 3300;
  localparam test_b1_S3301 = 3301;
  localparam test_b1_S3302 = 3302;
  localparam test_b1_S3303 = 3303;
  localparam test_b1_S3304 = 3304;
  localparam test_b1_S3305 = 3305;
  localparam test_b1_S3306 = 3306;
  localparam test_b1_S3307 = 3307;
  localparam test_b1_S3308 = 3308;
  localparam test_b1_S3309 = 3309;
  localparam test_b1_S3310 = 3310;
  localparam test_b1_S3311 = 3311;
  localparam test_b1_S3312 = 3312;
  localparam test_b1_S3313 = 3313;
  localparam test_b1_S3314 = 3314;
  localparam test_b1_S3315 = 3315;
  localparam test_b1_S3316 = 3316;
  localparam test_b1_S3317 = 3317;
  localparam test_b1_S3318 = 3318;
  localparam test_b1_S3319 = 3319;
  localparam test_b1_S3320 = 3320;
  localparam test_b1_S3321 = 3321;
  localparam test_b1_S3322 = 3322;
  localparam test_b1_S3323 = 3323;
  localparam test_b1_S3324 = 3324;
  localparam test_b1_S3325 = 3325;
  localparam test_b1_S3326 = 3326;
  localparam test_b1_S3327 = 3327;
  localparam test_b1_S3328 = 3328;
  localparam test_b1_S3329 = 3329;
  localparam test_b1_S3330 = 3330;
  localparam test_b1_S3331 = 3331;
  localparam test_b1_S3332 = 3332;
  localparam test_b1_S3333 = 3333;
  localparam test_b1_S3334 = 3334;
  localparam test_b1_S3335 = 3335;
  localparam test_b1_S3336 = 3336;
  localparam test_b1_S3337 = 3337;
  localparam test_b1_S3338 = 3338;
  localparam test_b1_S3339 = 3339;
  localparam test_b1_S3340 = 3340;
  localparam test_b1_S3341 = 3341;
  localparam test_b1_S3342 = 3342;
  localparam test_b1_S3343 = 3343;
  localparam test_b1_S3344 = 3344;
  localparam test_b1_S3345 = 3345;
  localparam test_b1_S3346 = 3346;
  localparam test_b1_S3347 = 3347;
  localparam test_b1_S3348 = 3348;
  localparam test_b1_S3349 = 3349;
  localparam test_b1_S3350 = 3350;
  localparam test_b1_S3351 = 3351;
  localparam test_b1_S3352 = 3352;
  localparam test_b1_S3353 = 3353;
  localparam test_b1_S3354 = 3354;
  localparam test_b1_S3355 = 3355;
  localparam test_b1_S3356 = 3356;
  localparam test_b1_S3357 = 3357;
  localparam test_b1_S3358 = 3358;
  localparam test_b1_S3359 = 3359;
  localparam test_b1_S3360 = 3360;
  localparam test_b1_S3361 = 3361;
  localparam test_b1_S3362 = 3362;
  localparam test_b1_S3363 = 3363;
  localparam test_b1_S3364 = 3364;
  localparam test_b1_S3365 = 3365;
  localparam test_b1_S3366 = 3366;
  localparam test_b1_S3367 = 3367;
  localparam test_b1_S3368 = 3368;
  localparam test_b1_S3369 = 3369;
  localparam test_b1_S3370 = 3370;
  localparam test_b1_S3371 = 3371;
  localparam test_b1_S3372 = 3372;
  localparam test_b1_S3373 = 3373;
  localparam test_b1_S3374 = 3374;
  localparam test_b1_S3375 = 3375;
  localparam test_b1_S3376 = 3376;
  localparam test_b1_S3377 = 3377;
  localparam test_b1_S3378 = 3378;
  localparam test_b1_S3379 = 3379;
  localparam test_b1_S3380 = 3380;
  localparam test_b1_S3381 = 3381;
  localparam test_b1_S3382 = 3382;
  localparam test_b1_S3383 = 3383;
  localparam test_b1_S3384 = 3384;
  localparam test_b1_S3385 = 3385;
  localparam test_b1_S3386 = 3386;
  localparam test_b1_S3387 = 3387;
  localparam test_b1_S3388 = 3388;
  localparam test_b1_S3389 = 3389;
  localparam test_b1_S3390 = 3390;
  localparam test_b1_S3391 = 3391;
  localparam test_b1_S3392 = 3392;
  localparam test_b1_S3393 = 3393;
  localparam test_b1_S3394 = 3394;
  localparam test_b1_S3395 = 3395;
  localparam test_b1_S3396 = 3396;
  localparam test_b1_S3397 = 3397;
  localparam test_b1_S3398 = 3398;
  localparam test_b1_S3399 = 3399;
  localparam test_b1_S3400 = 3400;
  localparam test_b1_S3401 = 3401;
  localparam test_b1_S3402 = 3402;
  localparam test_b1_S3403 = 3403;
  localparam test_b1_S3404 = 3404;
  localparam test_b1_S3405 = 3405;
  localparam test_b1_S3406 = 3406;
  localparam test_b1_S3407 = 3407;
  localparam test_b1_S3408 = 3408;
  localparam test_b1_S3409 = 3409;
  localparam test_b1_S3410 = 3410;
  localparam test_b1_S3411 = 3411;
  localparam test_b1_S3412 = 3412;
  localparam test_b1_S3413 = 3413;
  localparam test_b1_S3414 = 3414;
  localparam test_b1_S3415 = 3415;
  localparam test_b1_S3416 = 3416;
  localparam test_b1_S3417 = 3417;
  localparam test_b1_S3418 = 3418;
  localparam test_b1_S3419 = 3419;
  localparam test_b1_S3420 = 3420;
  localparam test_b1_S3421 = 3421;
  localparam test_b1_S3422 = 3422;
  localparam test_b1_S3423 = 3423;
  localparam test_b1_S3424 = 3424;
  localparam test_b1_S3425 = 3425;
  localparam test_b1_S3426 = 3426;
  localparam test_b1_S3427 = 3427;
  localparam test_b1_S3428 = 3428;
  localparam test_b1_S3429 = 3429;
  localparam test_b1_S3430 = 3430;
  localparam test_b1_S3431 = 3431;
  localparam test_b1_S3432 = 3432;
  localparam test_b1_S3433 = 3433;
  localparam test_b1_S3434 = 3434;
  localparam test_b1_S3435 = 3435;
  localparam test_b1_S3436 = 3436;
  localparam test_b1_S3437 = 3437;
  localparam test_b1_S3438 = 3438;
  localparam test_b1_S3439 = 3439;
  localparam test_b1_S3440 = 3440;
  localparam test_b1_S3441 = 3441;
  localparam test_b1_S3442 = 3442;
  localparam test_b1_S3443 = 3443;
  localparam test_b1_S3444 = 3444;
  localparam test_b1_S3445 = 3445;
  localparam test_b1_S3446 = 3446;
  localparam test_b1_S3447 = 3447;
  localparam test_b1_S3448 = 3448;
  localparam test_b1_S3449 = 3449;
  localparam test_b1_S3450 = 3450;
  localparam test_b1_S3451 = 3451;
  localparam test_b1_S3452 = 3452;
  localparam test_b1_S3453 = 3453;
  localparam test_b1_S3454 = 3454;
  localparam test_b1_S3455 = 3455;
  localparam test_b1_S3456 = 3456;
  localparam test_b1_S3457 = 3457;
  localparam test_b1_S3458 = 3458;
  localparam test_b1_S3459 = 3459;
  localparam test_b1_S3460 = 3460;
  localparam test_b1_S3461 = 3461;
  localparam test_b1_S3462 = 3462;
  localparam test_b1_S3463 = 3463;
  localparam test_b1_S3464 = 3464;
  localparam test_b1_S3465 = 3465;
  localparam test_b1_S3466 = 3466;
  localparam test_b1_S3467 = 3467;
  localparam test_b1_S3468 = 3468;
  localparam test_b1_S3469 = 3469;
  localparam test_b1_S3470 = 3470;
  localparam test_b1_S3471 = 3471;
  localparam test_b1_S3472 = 3472;
  localparam test_b1_S3473 = 3473;
  localparam test_b1_S3474 = 3474;
  localparam test_b1_S3475 = 3475;
  localparam test_b1_S3476 = 3476;
  localparam test_b1_S3477 = 3477;
  localparam test_b1_S3478 = 3478;
  localparam test_b1_S3479 = 3479;
  localparam test_b1_S3480 = 3480;
  localparam test_b1_S3481 = 3481;
  localparam test_b1_S3482 = 3482;
  localparam test_b1_S3483 = 3483;
  localparam test_b1_S3484 = 3484;
  localparam test_b1_S3485 = 3485;
  localparam test_b1_S3486 = 3486;
  localparam test_b1_S3487 = 3487;
  localparam test_b1_S3488 = 3488;
  localparam test_b1_S3489 = 3489;
  localparam test_b1_S3490 = 3490;
  localparam test_b1_S3491 = 3491;
  localparam test_b1_S3492 = 3492;
  localparam test_b1_S3493 = 3493;
  localparam test_b1_S3494 = 3494;
  localparam test_b1_S3495 = 3495;
  localparam test_b1_S3496 = 3496;
  localparam test_b1_S3497 = 3497;
  localparam test_b1_S3498 = 3498;
  localparam test_b1_S3499 = 3499;
  localparam test_b1_S3500 = 3500;
  localparam test_b1_S3501 = 3501;
  localparam test_b1_S3502 = 3502;
  localparam test_b1_S3503 = 3503;
  localparam test_b1_S3504 = 3504;
  localparam test_b1_S3505 = 3505;
  localparam test_b1_S3506 = 3506;
  localparam test_b1_S3507 = 3507;
  localparam test_b1_S3508 = 3508;
  localparam test_b1_S3509 = 3509;
  localparam test_b1_S3510 = 3510;
  localparam test_b1_S3511 = 3511;
  localparam test_b1_S3512 = 3512;
  localparam test_b1_S3513 = 3513;
  localparam test_b1_S3514 = 3514;
  localparam test_b1_S3515 = 3515;
  localparam test_b1_S3516 = 3516;
  localparam test_b1_S3517 = 3517;
  localparam test_b1_S3518 = 3518;
  localparam test_b1_S3519 = 3519;
  localparam test_b1_S3520 = 3520;
  localparam test_b1_S3521 = 3521;
  localparam test_b1_S3522 = 3522;
  localparam test_b1_S3523 = 3523;
  localparam test_b1_S3524 = 3524;
  localparam test_b1_S3525 = 3525;
  localparam test_b1_S3526 = 3526;
  localparam test_b1_S3527 = 3527;
  localparam test_b1_S3528 = 3528;
  localparam test_b1_S3529 = 3529;
  localparam test_b1_S3530 = 3530;
  localparam test_b1_S3531 = 3531;
  localparam test_b1_S3532 = 3532;
  localparam test_b1_S3533 = 3533;
  localparam test_b1_S3534 = 3534;
  localparam test_b1_S3535 = 3535;
  localparam test_b1_S3536 = 3536;
  localparam test_b1_S3537 = 3537;
  localparam test_b1_S3538 = 3538;
  localparam test_b1_S3539 = 3539;
  localparam test_b1_S3540 = 3540;
  localparam test_b1_S3541 = 3541;
  localparam test_b1_S3542 = 3542;
  localparam test_b1_S3543 = 3543;
  localparam test_b1_S3544 = 3544;
  localparam test_b1_S3545 = 3545;
  localparam test_b1_S3546 = 3546;
  localparam test_b1_S3547 = 3547;
  localparam test_b1_S3548 = 3548;
  localparam test_b1_S3549 = 3549;
  localparam test_b1_S3550 = 3550;
  localparam test_b1_S3551 = 3551;
  localparam test_b1_S3552 = 3552;
  localparam test_b1_S3553 = 3553;
  localparam test_b1_S3554 = 3554;
  localparam test_b1_S3555 = 3555;
  localparam test_b1_S3556 = 3556;
  localparam test_b1_S3557 = 3557;
  localparam test_b1_S3558 = 3558;
  localparam test_b1_S3559 = 3559;
  localparam test_b1_S3560 = 3560;
  localparam test_b1_S3561 = 3561;
  localparam test_b1_S3562 = 3562;
  localparam test_b1_S3563 = 3563;
  localparam test_b1_S3564 = 3564;
  localparam test_b1_S3565 = 3565;
  localparam test_b1_S3566 = 3566;
  localparam test_b1_S3567 = 3567;
  localparam test_b1_S3568 = 3568;
  localparam test_b1_S3569 = 3569;
  localparam test_b1_S3570 = 3570;
  localparam test_b1_S3571 = 3571;
  localparam test_b1_S3572 = 3572;
  localparam test_b1_S3573 = 3573;
  localparam test_b1_S3574 = 3574;
  localparam test_b1_S3575 = 3575;
  localparam test_b1_S3576 = 3576;
  localparam test_b1_S3577 = 3577;
  localparam test_b1_S3578 = 3578;
  localparam test_b1_S3579 = 3579;
  localparam test_b1_S3580 = 3580;
  localparam test_b1_S3581 = 3581;
  localparam test_b1_S3582 = 3582;
  localparam test_b1_S3583 = 3583;
  localparam test_b1_S3584 = 3584;
  localparam test_b1_S3585 = 3585;
  localparam test_b1_S3586 = 3586;
  localparam test_b1_S3587 = 3587;
  localparam test_b1_S3588 = 3588;
  localparam test_b1_S3589 = 3589;
  localparam test_b1_S3590 = 3590;
  localparam test_b1_S3591 = 3591;
  localparam test_b1_S3592 = 3592;
  localparam test_b1_S3593 = 3593;
  localparam test_b1_S3594 = 3594;
  localparam test_b1_S3595 = 3595;
  localparam test_b1_S3596 = 3596;
  localparam test_b1_S3597 = 3597;
  localparam test_b1_S3598 = 3598;
  localparam test_b1_S3599 = 3599;
  localparam test_b1_S3600 = 3600;
  localparam test_b1_S3601 = 3601;
  localparam test_b1_S3602 = 3602;
  localparam test_b1_S3603 = 3603;
  localparam test_b1_S3604 = 3604;
  localparam test_b1_S3605 = 3605;
  localparam test_b1_S3606 = 3606;
  localparam test_b1_S3607 = 3607;
  localparam test_b1_S3608 = 3608;
  localparam test_b1_S3609 = 3609;
  localparam test_b1_S3610 = 3610;
  localparam test_b1_S3611 = 3611;
  localparam test_b1_S3612 = 3612;
  localparam test_b1_S3613 = 3613;
  localparam test_b1_S3614 = 3614;
  localparam test_b1_S3615 = 3615;
  localparam test_b1_S3616 = 3616;
  localparam test_b1_S3617 = 3617;
  localparam test_b1_S3618 = 3618;
  localparam test_b1_S3619 = 3619;
  localparam test_b1_S3620 = 3620;
  localparam test_b1_S3621 = 3621;
  localparam test_b1_S3622 = 3622;
  localparam test_b1_S3623 = 3623;
  localparam test_b1_S3624 = 3624;
  localparam test_b1_S3625 = 3625;
  localparam test_b1_S3626 = 3626;
  localparam test_b1_S3627 = 3627;
  localparam test_b1_S3628 = 3628;
  localparam test_b1_S3629 = 3629;
  localparam test_b1_S3630 = 3630;
  localparam test_b1_S3631 = 3631;
  localparam test_b1_S3632 = 3632;
  localparam test_b1_S3633 = 3633;
  localparam test_b1_S3634 = 3634;
  localparam test_b1_S3635 = 3635;
  localparam test_b1_S3636 = 3636;
  localparam test_b1_S3637 = 3637;
  localparam test_b1_S3638 = 3638;
  localparam test_b1_S3639 = 3639;
  localparam test_b1_S3640 = 3640;
  localparam test_b1_S3641 = 3641;
  localparam test_b1_S3642 = 3642;
  localparam test_b1_S3643 = 3643;
  localparam test_b1_S3644 = 3644;
  localparam test_b1_S3645 = 3645;
  localparam test_b1_S3646 = 3646;
  localparam test_b1_S3647 = 3647;
  localparam test_b1_S3648 = 3648;
  localparam test_b1_S3649 = 3649;
  localparam test_b1_S3650 = 3650;
  localparam test_b1_S3651 = 3651;
  localparam test_b1_S3652 = 3652;
  localparam test_b1_S3653 = 3653;
  localparam test_b1_S3654 = 3654;
  localparam test_b1_S3655 = 3655;
  localparam test_b1_S3656 = 3656;
  localparam test_b1_S3657 = 3657;
  localparam test_b1_S3658 = 3658;
  localparam test_b1_S3659 = 3659;
  localparam test_b1_S3660 = 3660;
  localparam test_b1_S3661 = 3661;
  localparam test_b1_S3662 = 3662;
  localparam test_b1_S3663 = 3663;
  localparam test_b1_S3664 = 3664;
  localparam test_b1_S3665 = 3665;
  localparam test_b1_S3666 = 3666;
  localparam test_b1_S3667 = 3667;
  localparam test_b1_S3668 = 3668;
  localparam test_b1_S3669 = 3669;
  localparam test_b1_S3670 = 3670;
  localparam test_b1_S3671 = 3671;
  localparam test_b1_S3672 = 3672;
  localparam test_b1_S3673 = 3673;
  localparam test_b1_S3674 = 3674;
  localparam test_b1_S3675 = 3675;
  localparam test_b1_S3676 = 3676;
  localparam test_b1_S3677 = 3677;
  localparam test_b1_S3678 = 3678;
  localparam test_b1_S3679 = 3679;
  localparam test_b1_S3680 = 3680;
  localparam test_b1_S3681 = 3681;
  localparam test_b1_S3682 = 3682;
  localparam test_b1_S3683 = 3683;
  localparam test_b1_S3684 = 3684;
  localparam test_b1_S3685 = 3685;
  localparam test_b1_S3686 = 3686;
  localparam test_b1_S3687 = 3687;
  localparam test_b1_S3688 = 3688;
  localparam test_b1_S3689 = 3689;
  localparam test_b1_S3690 = 3690;
  localparam test_b1_S3691 = 3691;
  localparam test_b1_S3692 = 3692;
  localparam test_b1_S3693 = 3693;
  localparam test_b1_S3694 = 3694;
  localparam test_b1_S3695 = 3695;
  localparam test_b1_S3696 = 3696;
  localparam test_b1_S3697 = 3697;
  localparam test_b1_S3698 = 3698;
  localparam test_b1_S3699 = 3699;
  localparam test_b1_S3700 = 3700;
  localparam test_b1_S3701 = 3701;
  localparam test_b1_S3702 = 3702;
  localparam test_b1_S3703 = 3703;
  localparam test_b1_S3704 = 3704;
  localparam test_b1_S3705 = 3705;
  localparam test_b1_S3706 = 3706;
  localparam test_b1_S3707 = 3707;
  localparam test_b1_S3708 = 3708;
  localparam test_b1_S3709 = 3709;
  localparam test_b1_S3710 = 3710;
  localparam test_b1_S3711 = 3711;
  localparam test_b1_S3712 = 3712;
  localparam test_b1_S3713 = 3713;
  localparam test_b1_S3714 = 3714;
  localparam test_b1_S3715 = 3715;
  localparam test_b1_S3716 = 3716;
  localparam test_b1_S3717 = 3717;
  localparam test_b1_S3718 = 3718;
  localparam test_b1_S3719 = 3719;
  localparam test_b1_S3720 = 3720;
  localparam test_b1_S3721 = 3721;
  localparam test_b1_S3722 = 3722;
  localparam test_b1_S3723 = 3723;
  localparam test_b1_S3724 = 3724;
  localparam test_b1_S3725 = 3725;
  localparam test_b1_S3726 = 3726;
  localparam test_b1_S3727 = 3727;
  localparam test_b1_S3728 = 3728;
  localparam test_b1_S3729 = 3729;
  localparam test_b1_S3730 = 3730;
  localparam test_b1_S3731 = 3731;
  localparam test_b1_S3732 = 3732;
  localparam test_b1_S3733 = 3733;
  localparam test_b1_S3734 = 3734;
  localparam test_b1_S3735 = 3735;
  localparam test_b1_S3736 = 3736;
  localparam test_b1_S3737 = 3737;
  localparam test_b1_S3738 = 3738;
  localparam test_b1_S3739 = 3739;
  localparam test_b1_S3740 = 3740;
  localparam test_b1_S3741 = 3741;
  localparam test_b1_S3742 = 3742;
  localparam test_b1_S3743 = 3743;
  localparam test_b1_S3744 = 3744;
  localparam test_b1_S3745 = 3745;
  localparam test_b1_S3746 = 3746;
  localparam test_b1_S3747 = 3747;
  localparam test_b1_S3748 = 3748;
  localparam test_b1_S3749 = 3749;
  localparam test_b1_S3750 = 3750;
  localparam test_b1_S3751 = 3751;
  localparam test_b1_S3752 = 3752;
  localparam test_b1_S3753 = 3753;
  localparam test_b1_S3754 = 3754;
  localparam test_b1_S3755 = 3755;
  localparam test_b1_S3756 = 3756;
  localparam test_b1_S3757 = 3757;
  localparam test_b1_S3758 = 3758;
  localparam test_b1_S3759 = 3759;
  localparam test_b1_S3760 = 3760;
  localparam test_b1_S3761 = 3761;
  localparam test_b1_S3762 = 3762;
  localparam test_b1_S3763 = 3763;
  localparam test_b1_S3764 = 3764;
  localparam test_b1_S3765 = 3765;
  localparam test_b1_S3766 = 3766;
  localparam test_b1_S3767 = 3767;
  localparam test_b1_S3768 = 3768;
  localparam test_b1_S3769 = 3769;
  localparam test_b1_S3770 = 3770;
  localparam test_b1_S3771 = 3771;
  localparam test_b1_S3772 = 3772;
  localparam test_b1_S3773 = 3773;
  localparam test_b1_S3774 = 3774;
  localparam test_b1_S3775 = 3775;
  localparam test_b1_S3776 = 3776;
  localparam test_b1_S3777 = 3777;
  localparam test_b1_S3778 = 3778;
  localparam test_b1_S3779 = 3779;
  localparam test_b1_S3780 = 3780;
  localparam test_b1_S3781 = 3781;
  localparam test_b1_S3782 = 3782;
  localparam test_b1_S3783 = 3783;
  localparam test_b1_S3784 = 3784;
  localparam test_b1_S3785 = 3785;
  localparam test_b1_S3786 = 3786;
  localparam test_b1_S3787 = 3787;
  localparam test_b1_S3788 = 3788;
  localparam test_b1_S3789 = 3789;
  localparam test_b1_S3790 = 3790;
  localparam test_b1_S3791 = 3791;
  localparam test_b1_S3792 = 3792;
  localparam test_b1_S3793 = 3793;
  localparam test_b1_S3794 = 3794;
  localparam test_b1_S3795 = 3795;
  localparam test_b1_S3796 = 3796;
  localparam test_b1_S3797 = 3797;
  localparam test_b1_S3798 = 3798;
  localparam test_b1_S3799 = 3799;
  localparam test_b1_S3800 = 3800;
  localparam test_b1_S3801 = 3801;
  localparam test_b1_S3802 = 3802;
  localparam test_b1_S3803 = 3803;
  localparam test_b1_S3804 = 3804;
  localparam test_b1_S3805 = 3805;
  localparam test_b1_S3806 = 3806;
  localparam test_b1_S3807 = 3807;
  localparam test_b1_S3808 = 3808;
  localparam test_b1_S3809 = 3809;
  localparam test_b1_S3810 = 3810;
  localparam test_b1_S3811 = 3811;
  localparam test_b1_S3812 = 3812;
  localparam test_b1_S3813 = 3813;
  localparam test_b1_S3814 = 3814;
  localparam test_b1_S3815 = 3815;
  localparam test_b1_S3816 = 3816;
  localparam test_b1_S3817 = 3817;
  localparam test_b1_S3818 = 3818;
  localparam test_b1_S3819 = 3819;
  localparam test_b1_S3820 = 3820;
  localparam test_b1_S3821 = 3821;
  localparam test_b1_S3822 = 3822;
  localparam test_b1_S3823 = 3823;
  localparam test_b1_S3824 = 3824;
  localparam test_b1_S3825 = 3825;
  localparam test_b1_S3826 = 3826;
  localparam test_b1_S3827 = 3827;
  localparam test_b1_S3828 = 3828;
  localparam test_b1_S3829 = 3829;
  localparam test_b1_S3830 = 3830;
  localparam test_b1_S3831 = 3831;
  localparam test_b1_S3832 = 3832;
  localparam test_b1_S3833 = 3833;
  localparam test_b1_S3834 = 3834;
  localparam test_b1_S3835 = 3835;
  localparam test_b1_S3836 = 3836;
  localparam test_b1_S3837 = 3837;
  localparam test_b1_S3838 = 3838;
  localparam test_b1_S3839 = 3839;
  localparam test_b1_S3840 = 3840;
  localparam test_b1_S3841 = 3841;
  localparam test_b1_S3842 = 3842;
  localparam test_b1_S3843 = 3843;
  localparam test_b1_S3844 = 3844;
  localparam test_b1_S3845 = 3845;
  localparam test_b1_S3846 = 3846;
  localparam test_b1_S3847 = 3847;
  localparam test_b1_S3848 = 3848;
  localparam test_b1_S3849 = 3849;
  localparam test_b1_S3850 = 3850;
  localparam test_b1_S3851 = 3851;
  localparam test_b1_S3852 = 3852;
  localparam test_b1_S3853 = 3853;
  localparam test_b1_S3854 = 3854;
  localparam test_b1_S3855 = 3855;
  localparam test_b1_S3856 = 3856;
  localparam test_b1_S3857 = 3857;
  localparam test_b1_S3858 = 3858;
  localparam test_b1_S3859 = 3859;
  localparam test_b1_S3860 = 3860;
  localparam test_b1_S3861 = 3861;
  localparam test_b1_S3862 = 3862;
  localparam test_b1_S3863 = 3863;
  localparam test_b1_S3864 = 3864;
  localparam test_b1_S3865 = 3865;
  localparam test_b1_S3866 = 3866;
  localparam test_b1_S3867 = 3867;
  localparam test_b1_S3868 = 3868;
  localparam test_b1_S3869 = 3869;
  localparam test_b1_S3870 = 3870;
  localparam test_b1_S3871 = 3871;
  localparam test_b1_S3872 = 3872;
  localparam test_b1_S3873 = 3873;
  localparam test_b1_S3874 = 3874;
  localparam test_b1_S3875 = 3875;
  localparam test_b1_S3876 = 3876;
  localparam test_b1_S3877 = 3877;
  localparam test_b1_S3878 = 3878;
  localparam test_b1_S3879 = 3879;
  localparam test_b1_S3880 = 3880;
  localparam test_b1_S3881 = 3881;
  localparam test_b1_S3882 = 3882;
  localparam test_b1_S3883 = 3883;
  localparam test_b1_S3884 = 3884;
  localparam test_b1_S3885 = 3885;
  localparam test_b1_S3886 = 3886;
  localparam test_b1_S3887 = 3887;
  localparam test_b1_S3888 = 3888;
  localparam test_b1_S3889 = 3889;
  localparam test_b1_S3890 = 3890;
  localparam test_b1_S3891 = 3891;
  localparam test_b1_S3892 = 3892;
  localparam test_b1_S3893 = 3893;
  localparam test_b1_S3894 = 3894;
  localparam test_b1_S3895 = 3895;
  localparam test_b1_S3896 = 3896;
  localparam test_b1_S3897 = 3897;
  localparam test_b1_S3898 = 3898;
  localparam test_b1_S3899 = 3899;
  localparam test_b1_S3900 = 3900;
  localparam test_b1_S3901 = 3901;
  localparam test_b1_S3902 = 3902;
  localparam test_b1_S3903 = 3903;
  localparam test_b1_S3904 = 3904;
  localparam test_b1_S3905 = 3905;
  localparam test_b1_S3906 = 3906;
  localparam test_b1_S3907 = 3907;
  localparam test_b1_S3908 = 3908;
  localparam test_b1_S3909 = 3909;
  localparam test_b1_S3910 = 3910;
  localparam test_b1_S3911 = 3911;
  localparam test_b1_S3912 = 3912;
  localparam test_b1_S3913 = 3913;
  localparam test_b1_S3914 = 3914;
  localparam test_b1_S3915 = 3915;
  localparam test_b1_S3916 = 3916;
  localparam test_b1_S3917 = 3917;
  localparam test_b1_S3918 = 3918;
  localparam test_b1_S3919 = 3919;
  localparam test_b1_S3920 = 3920;
  localparam test_b1_S3921 = 3921;
  localparam test_b1_S3922 = 3922;
  localparam test_b1_S3923 = 3923;
  localparam test_b1_S3924 = 3924;
  localparam test_b1_S3925 = 3925;
  localparam test_b1_S3926 = 3926;
  localparam test_b1_S3927 = 3927;
  localparam test_b1_S3928 = 3928;
  localparam test_b1_S3929 = 3929;
  localparam test_b1_S3930 = 3930;
  localparam test_b1_S3931 = 3931;
  localparam test_b1_S3932 = 3932;
  localparam test_b1_S3933 = 3933;
  localparam test_b1_S3934 = 3934;
  localparam test_b1_S3935 = 3935;
  localparam test_b1_S3936 = 3936;
  localparam test_b1_S3937 = 3937;
  localparam test_b1_S3938 = 3938;
  localparam test_b1_S3939 = 3939;
  localparam test_b1_S3940 = 3940;
  localparam test_b1_S3941 = 3941;
  localparam test_b1_S3942 = 3942;
  localparam test_b1_S3943 = 3943;
  localparam test_b1_S3944 = 3944;
  localparam test_b1_S3945 = 3945;
  localparam test_b1_S3946 = 3946;
  localparam test_b1_S3947 = 3947;
  localparam test_b1_S3948 = 3948;
  localparam test_b1_S3949 = 3949;
  localparam test_b1_S3950 = 3950;
  localparam test_b1_S3951 = 3951;
  localparam test_b1_S3952 = 3952;
  localparam test_b1_S3953 = 3953;
  localparam test_b1_S3954 = 3954;
  localparam test_b1_S3955 = 3955;
  localparam test_b1_S3956 = 3956;
  localparam test_b1_S3957 = 3957;
  localparam test_b1_S3958 = 3958;
  localparam test_b1_S3959 = 3959;
  localparam test_b1_S3960 = 3960;
  localparam test_b1_S3961 = 3961;
  localparam test_b1_S3962 = 3962;
  localparam test_b1_S3963 = 3963;
  localparam test_b1_S3964 = 3964;
  localparam test_b1_S3965 = 3965;
  localparam test_b1_S3966 = 3966;
  localparam test_b1_S3967 = 3967;
  localparam test_b1_S3968 = 3968;
  localparam test_b1_S3969 = 3969;
  localparam test_b1_S3970 = 3970;
  localparam test_b1_S3971 = 3971;
  localparam test_b1_S3972 = 3972;
  localparam test_b1_S3973 = 3973;
  localparam test_b1_S3974 = 3974;
  localparam test_b1_S3975 = 3975;
  localparam test_b1_S3976 = 3976;
  localparam test_b1_S3977 = 3977;
  localparam test_b1_S3978 = 3978;
  localparam test_b1_S3979 = 3979;
  localparam test_b1_S3980 = 3980;
  localparam test_b1_S3981 = 3981;
  localparam test_b1_S3982 = 3982;
  localparam test_b1_S3983 = 3983;
  localparam test_b1_S3984 = 3984;
  localparam test_b1_S3985 = 3985;
  localparam test_b1_S3986 = 3986;
  localparam test_b1_S3987 = 3987;
  localparam test_b1_S3988 = 3988;
  localparam test_b1_S3989 = 3989;
  localparam test_b1_S3990 = 3990;
  localparam test_b1_S3991 = 3991;
  localparam test_b1_S3992 = 3992;
  localparam test_b1_S3993 = 3993;
  localparam test_b1_S3994 = 3994;
  localparam test_b1_S3995 = 3995;
  localparam test_b1_S3996 = 3996;
  localparam test_b1_S3997 = 3997;
  localparam test_b1_S3998 = 3998;
  localparam test_b1_S3999 = 3999;
  localparam test_b1_S4000 = 4000;
  localparam test_b1_S4001 = 4001;
  localparam test_b1_S4002 = 4002;
  localparam test_b1_S4003 = 4003;
  localparam test_b1_S4004 = 4004;
  localparam test_b1_S4005 = 4005;
  localparam test_b1_S4006 = 4006;
  localparam test_b1_S4007 = 4007;
  localparam test_b1_S4008 = 4008;
  localparam test_b1_S4009 = 4009;
  localparam test_b1_S4010 = 4010;
  localparam test_b1_S4011 = 4011;
  localparam test_b1_S4012 = 4012;
  localparam test_b1_S4013 = 4013;
  localparam test_b1_S4014 = 4014;
  localparam test_b1_S4015 = 4015;
  localparam test_b1_S4016 = 4016;
  localparam test_b1_S4017 = 4017;
  localparam test_b1_S4018 = 4018;
  localparam test_b1_S4019 = 4019;
  localparam test_b1_S4020 = 4020;
  localparam test_b1_S4021 = 4021;
  localparam test_b1_S4022 = 4022;
  localparam test_b1_S4023 = 4023;
  localparam test_b1_S4024 = 4024;
  localparam test_b1_S4025 = 4025;
  localparam test_b1_S4026 = 4026;
  localparam test_b1_S4027 = 4027;
  localparam test_b1_S4028 = 4028;
  localparam test_b1_S4029 = 4029;
  localparam test_b1_S4030 = 4030;
  localparam test_b1_S4031 = 4031;
  localparam test_b1_S4032 = 4032;
  localparam test_b1_S4033 = 4033;
  localparam test_b1_S4034 = 4034;
  localparam test_b1_S4035 = 4035;
  localparam test_b1_S4036 = 4036;
  localparam test_b1_S4037 = 4037;
  localparam test_b1_S4038 = 4038;
  localparam test_b1_S4039 = 4039;
  localparam test_b1_S4040 = 4040;
  localparam test_b1_S4041 = 4041;
  localparam test_b1_S4042 = 4042;
  localparam test_b1_S4043 = 4043;
  localparam test_b1_S4044 = 4044;
  localparam test_b1_S4045 = 4045;
  localparam test_b1_S4046 = 4046;
  localparam test_b1_S4047 = 4047;
  localparam test_b1_S4048 = 4048;
  localparam test_b1_S4049 = 4049;
  localparam test_b1_S4050 = 4050;
  localparam test_b1_S4051 = 4051;
  localparam test_b1_S4052 = 4052;
  localparam test_b1_S4053 = 4053;
  localparam test_b1_S4054 = 4054;
  localparam test_b1_S4055 = 4055;
  localparam test_b1_S4056 = 4056;
  localparam test_b1_S4057 = 4057;
  localparam test_b1_S4058 = 4058;
  localparam test_b1_S4059 = 4059;
  localparam test_b1_S4060 = 4060;
  localparam test_b1_S4061 = 4061;
  localparam test_b1_S4062 = 4062;
  localparam test_b1_S4063 = 4063;
  localparam test_b1_S4064 = 4064;
  localparam test_b1_S4065 = 4065;
  localparam test_b1_S4066 = 4066;
  localparam test_b1_S4067 = 4067;
  localparam test_b1_S4068 = 4068;
  localparam test_b1_S4069 = 4069;
  localparam test_b1_S4070 = 4070;
  localparam test_b1_S4071 = 4071;
  localparam test_b1_S4072 = 4072;
  localparam test_b1_S4073 = 4073;
  localparam test_b1_S4074 = 4074;
  localparam test_b1_S4075 = 4075;
  localparam test_b1_S4076 = 4076;
  localparam test_b1_S4077 = 4077;
  localparam test_b1_S4078 = 4078;
  localparam test_b1_S4079 = 4079;
  localparam test_b1_S4080 = 4080;
  localparam test_b1_S4081 = 4081;
  localparam test_b1_S4082 = 4082;
  localparam test_b1_S4083 = 4083;
  localparam test_b1_S4084 = 4084;
  localparam test_b1_S4085 = 4085;
  localparam test_b1_S4086 = 4086;
  localparam test_b1_S4087 = 4087;
  localparam test_b1_S4088 = 4088;
  localparam test_b1_S4089 = 4089;
  localparam test_b1_S4090 = 4090;
  localparam test_b1_S4091 = 4091;
  localparam test_b1_S4092 = 4092;
  localparam test_b1_S4093 = 4093;
  localparam test_b1_S4094 = 4094;
  localparam test_b1_S4095 = 4095;
  localparam test_b1_S4096 = 4096;
  localparam test_b1_S4097 = 4097;
  localparam test_b1_S4098 = 4098;
  localparam test_b1_S4099 = 4099;
  localparam test_b1_S4100 = 4100;
  localparam test_b1_S4101 = 4101;
  localparam test_b1_S4102 = 4102;
  localparam test_b1_S4103 = 4103;
  localparam test_b1_S4104 = 4104;
  localparam test_b1_S4105 = 4105;
  localparam test_b1_S4106 = 4106;
  localparam test_b1_S4107 = 4107;
  localparam test_b1_S4108 = 4108;
  localparam test_b1_S4109 = 4109;
  localparam test_b1_S4110 = 4110;
  localparam test_b1_S4111 = 4111;
  localparam test_b1_S4112 = 4112;
  localparam test_b1_S4113 = 4113;
  localparam test_b1_S4114 = 4114;
  localparam test_b1_S4115 = 4115;
  localparam test_b1_S4116 = 4116;
  localparam test_b1_S4117 = 4117;
  localparam test_b1_S4118 = 4118;
  localparam test_b1_S4119 = 4119;
  localparam test_b1_S4120 = 4120;
  localparam test_b1_S4121 = 4121;
  localparam test_b1_S4122 = 4122;
  localparam test_b1_S4123 = 4123;
  localparam test_b1_S4124 = 4124;
  localparam test_b1_S4125 = 4125;
  localparam test_b1_S4126 = 4126;
  localparam test_b1_S4127 = 4127;
  localparam test_b1_S4128 = 4128;
  localparam test_b1_S4129 = 4129;
  localparam test_b1_S4130 = 4130;
  localparam test_b1_S4131 = 4131;
  localparam test_b1_S4132 = 4132;
  localparam test_b1_S4133 = 4133;
  localparam test_b1_S4134 = 4134;
  localparam test_b1_S4135 = 4135;
  localparam test_b1_S4136 = 4136;
  localparam test_b1_S4137 = 4137;
  localparam test_b1_S4138 = 4138;
  localparam test_b1_S4139 = 4139;
  localparam test_b1_S4140 = 4140;
  localparam test_b1_S4141 = 4141;
  localparam test_b1_S4142 = 4142;
  localparam test_b1_S4143 = 4143;
  localparam test_b1_S4144 = 4144;
  localparam test_b1_S4145 = 4145;
  localparam test_b1_S4146 = 4146;
  localparam test_b1_S4147 = 4147;
  localparam test_b1_S4148 = 4148;
  localparam test_b1_S4149 = 4149;
  localparam test_b1_S4150 = 4150;
  localparam test_b1_S4151 = 4151;
  localparam test_b1_S4152 = 4152;
  localparam test_b1_S4153 = 4153;
  localparam test_b1_S4154 = 4154;
  localparam test_b1_S4155 = 4155;
  localparam test_b1_S4156 = 4156;
  localparam test_b1_S4157 = 4157;
  localparam test_b1_S4158 = 4158;
  localparam test_b1_S4159 = 4159;
  localparam test_b1_S4160 = 4160;
  localparam test_b1_S4161 = 4161;
  localparam test_b1_S4162 = 4162;
  localparam test_b1_S4163 = 4163;
  localparam test_b1_S4164 = 4164;
  localparam test_b1_S4165 = 4165;
  localparam test_b1_S4166 = 4166;
  localparam test_b1_S4167 = 4167;
  localparam test_b1_S4168 = 4168;
  localparam test_b1_S4169 = 4169;
  localparam test_b1_S4170 = 4170;
  localparam test_b1_S4171 = 4171;
  localparam test_b1_S4172 = 4172;
  localparam test_b1_S4173 = 4173;
  localparam test_b1_S4174 = 4174;
  localparam test_b1_S4175 = 4175;
  localparam test_b1_S4176 = 4176;
  localparam test_b1_S4177 = 4177;
  localparam test_b1_S4178 = 4178;
  localparam test_b1_S4179 = 4179;
  localparam test_b1_S4180 = 4180;
  localparam test_b1_S4181 = 4181;
  localparam test_b1_S4182 = 4182;
  localparam test_b1_S4183 = 4183;
  localparam test_b1_S4184 = 4184;
  localparam test_b1_S4185 = 4185;
  localparam test_b1_S4186 = 4186;
  localparam test_b1_S4187 = 4187;
  localparam test_b1_S4188 = 4188;
  localparam test_b1_S4189 = 4189;
  localparam test_b1_S4190 = 4190;
  localparam test_b1_S4191 = 4191;
  localparam test_b1_S4192 = 4192;
  localparam test_b1_S4193 = 4193;
  localparam test_b1_S4194 = 4194;
  localparam test_b1_S4195 = 4195;
  localparam test_b1_S4196 = 4196;
  localparam test_b1_S4197 = 4197;
  localparam test_b1_S4198 = 4198;
  localparam test_b1_S4199 = 4199;
  localparam test_b1_S4200 = 4200;
  localparam test_b1_S4201 = 4201;
  localparam test_b1_S4202 = 4202;
  localparam test_b1_S4203 = 4203;
  localparam test_b1_S4204 = 4204;
  localparam test_b1_S4205 = 4205;
  localparam test_b1_S4206 = 4206;
  localparam test_b1_S4207 = 4207;
  localparam test_b1_S4208 = 4208;
  localparam test_b1_S4209 = 4209;
  localparam test_b1_S4210 = 4210;
  localparam test_b1_S4211 = 4211;
  localparam test_b1_S4212 = 4212;
  localparam test_b1_S4213 = 4213;
  localparam test_b1_S4214 = 4214;
  localparam test_b1_S4215 = 4215;
  localparam test_b1_S4216 = 4216;
  localparam test_b1_S4217 = 4217;
  localparam test_b1_S4218 = 4218;
  localparam test_b1_S4219 = 4219;
  localparam test_b1_S4220 = 4220;
  localparam test_b1_S4221 = 4221;
  localparam test_b1_S4222 = 4222;
  localparam test_b1_S4223 = 4223;
  localparam test_b1_S4224 = 4224;
  localparam test_b1_S4225 = 4225;
  localparam test_b1_S4226 = 4226;
  localparam test_b1_S4227 = 4227;
  localparam test_b1_S4228 = 4228;
  localparam test_b1_S4229 = 4229;
  localparam test_b1_S4230 = 4230;
  localparam test_b1_S4231 = 4231;
  localparam test_b1_S4232 = 4232;
  localparam test_b1_S4233 = 4233;
  localparam test_b1_S4234 = 4234;
  localparam test_b1_S4235 = 4235;
  localparam test_b1_S4236 = 4236;
  localparam test_b1_S4237 = 4237;
  localparam test_b1_S4238 = 4238;
  localparam test_b1_S4239 = 4239;
  localparam test_b1_S4240 = 4240;
  localparam test_b1_S4241 = 4241;
  localparam test_b1_S4242 = 4242;
  localparam test_b1_S4243 = 4243;
  localparam test_b1_S4244 = 4244;
  localparam test_b1_S4245 = 4245;
  localparam test_b1_S4246 = 4246;
  localparam test_b1_S4247 = 4247;
  localparam test_b1_S4248 = 4248;
  localparam test_b1_S4249 = 4249;
  localparam test_b1_S4250 = 4250;
  localparam test_b1_S4251 = 4251;
  localparam test_b1_S4252 = 4252;
  localparam test_b1_S4253 = 4253;
  localparam test_b1_S4254 = 4254;
  localparam test_b1_S4255 = 4255;
  localparam test_b1_S4256 = 4256;
  localparam test_b1_S4257 = 4257;
  localparam test_b1_S4258 = 4258;
  localparam test_b1_S4259 = 4259;
  localparam test_b1_S4260 = 4260;
  localparam test_b1_S4261 = 4261;
  localparam test_b1_S4262 = 4262;
  localparam test_b1_S4263 = 4263;
  localparam test_b1_S4264 = 4264;
  localparam test_b1_S4265 = 4265;
  localparam test_b1_S4266 = 4266;
  localparam test_b1_S4267 = 4267;
  localparam test_b1_S4268 = 4268;
  localparam test_b1_S4269 = 4269;
  localparam test_b1_S4270 = 4270;
  localparam test_b1_S4271 = 4271;
  localparam test_b1_S4272 = 4272;
  localparam test_b1_S4273 = 4273;
  localparam test_b1_S4274 = 4274;
  localparam test_b1_S4275 = 4275;
  localparam test_b1_S4276 = 4276;
  localparam test_b1_S4277 = 4277;
  localparam test_b1_S4278 = 4278;
  localparam test_b1_S4279 = 4279;
  localparam test_b1_S4280 = 4280;
  localparam test_b1_S4281 = 4281;
  localparam test_b1_S4282 = 4282;
  localparam test_b1_S4283 = 4283;
  localparam test_b1_S4284 = 4284;
  localparam test_b1_S4285 = 4285;
  localparam test_b1_S4286 = 4286;
  localparam test_b1_S4287 = 4287;
  localparam test_b1_S4288 = 4288;
  localparam test_b1_S4289 = 4289;
  localparam test_b1_S4290 = 4290;
  localparam test_b1_S4291 = 4291;
  localparam test_b1_S4292 = 4292;
  localparam test_b1_S4293 = 4293;
  localparam test_b1_S4294 = 4294;
  localparam test_b1_S4295 = 4295;
  localparam test_b1_S4296 = 4296;
  localparam test_b1_S4297 = 4297;
  localparam test_b1_S4298 = 4298;
  localparam test_b1_S4299 = 4299;
  localparam test_b1_S4300 = 4300;
  localparam test_b1_S4301 = 4301;
  localparam test_b1_S4302 = 4302;
  localparam test_b1_S4303 = 4303;
  localparam test_b1_S4304 = 4304;
  localparam test_b1_S4305 = 4305;
  localparam test_b1_S4306 = 4306;
  localparam test_b1_S4307 = 4307;
  localparam test_b1_S4308 = 4308;
  localparam test_b1_S4309 = 4309;
  localparam test_b1_S4310 = 4310;
  localparam test_b1_S4311 = 4311;
  localparam test_b1_S4312 = 4312;
  localparam test_b1_S4313 = 4313;
  localparam test_b1_S4314 = 4314;
  localparam test_b1_S4315 = 4315;
  localparam test_b1_S4316 = 4316;
  localparam test_b1_S4317 = 4317;
  localparam test_b1_S4318 = 4318;
  localparam test_b1_S4319 = 4319;
  localparam test_b1_S4320 = 4320;
  localparam test_b1_S4321 = 4321;
  localparam test_b1_S4322 = 4322;
  localparam test_b1_S4323 = 4323;
  localparam test_b1_S4324 = 4324;
  localparam test_b1_S4325 = 4325;
  localparam test_b1_S4326 = 4326;
  localparam test_b1_S4327 = 4327;
  localparam test_b1_S4328 = 4328;
  localparam test_b1_S4329 = 4329;
  localparam test_b1_S4330 = 4330;
  localparam test_b1_S4331 = 4331;
  localparam test_b1_S4332 = 4332;
  localparam test_b1_S4333 = 4333;
  localparam test_b1_S4334 = 4334;
  localparam test_b1_S4335 = 4335;
  localparam test_b1_S4336 = 4336;
  localparam test_b1_S4337 = 4337;
  localparam test_b1_S4338 = 4338;
  localparam test_b1_S4339 = 4339;
  localparam test_b1_S4340 = 4340;
  localparam test_b1_S4341 = 4341;
  localparam test_b1_S4342 = 4342;
  localparam test_b1_S4343 = 4343;
  localparam test_b1_S4344 = 4344;
  localparam test_b1_S4345 = 4345;
  localparam test_b1_S4346 = 4346;
  localparam test_b1_S4347 = 4347;
  localparam test_b1_S4348 = 4348;
  localparam test_b1_S4349 = 4349;
  localparam test_b1_S4350 = 4350;
  localparam test_b1_S4351 = 4351;
  localparam test_b1_S4352 = 4352;
  localparam test_b1_S4353 = 4353;
  localparam test_b1_S4354 = 4354;
  localparam test_b1_S4355 = 4355;
  localparam test_b1_S4356 = 4356;
  localparam test_b1_S4357 = 4357;
  localparam test_b1_S4358 = 4358;
  localparam test_b1_S4359 = 4359;
  localparam test_b1_S4360 = 4360;
  localparam test_b1_S4361 = 4361;
  localparam test_b1_S4362 = 4362;
  localparam test_b1_S4363 = 4363;
  localparam test_b1_S4364 = 4364;
  localparam test_b1_S4365 = 4365;
  localparam test_b1_S4366 = 4366;
  localparam test_b1_S4367 = 4367;
  localparam test_b1_S4368 = 4368;
  localparam test_b1_S4369 = 4369;
  localparam test_b1_S4370 = 4370;
  localparam test_b1_S4371 = 4371;
  localparam test_b1_S4372 = 4372;
  localparam test_b1_S4373 = 4373;
  localparam test_b1_S4374 = 4374;
  localparam test_b1_S4375 = 4375;
  localparam test_b1_S4376 = 4376;
  localparam test_b1_S4377 = 4377;
  localparam test_b1_S4378 = 4378;
  localparam test_b1_S4379 = 4379;
  localparam test_b1_S4380 = 4380;
  localparam test_b1_S4381 = 4381;
  localparam test_b1_S4382 = 4382;
  localparam test_b1_S4383 = 4383;
  localparam test_b1_S4384 = 4384;
  localparam test_b1_S4385 = 4385;
  localparam test_b1_S4386 = 4386;
  localparam test_b1_S4387 = 4387;
  localparam test_b1_S4388 = 4388;
  localparam test_b1_S4389 = 4389;
  localparam test_b1_S4390 = 4390;
  localparam test_b1_S4391 = 4391;
  localparam test_b1_S4392 = 4392;
  localparam test_b1_S4393 = 4393;
  localparam test_b1_S4394 = 4394;
  localparam test_b1_S4395 = 4395;
  localparam test_b1_S4396 = 4396;
  localparam test_b1_S4397 = 4397;
  localparam test_b1_S4398 = 4398;
  localparam test_b1_S4399 = 4399;
  localparam test_b1_S4400 = 4400;
  localparam test_b1_S4401 = 4401;
  localparam test_b1_S4402 = 4402;
  localparam test_b1_S4403 = 4403;
  localparam test_b1_S4404 = 4404;
  localparam test_b1_S4405 = 4405;
  localparam test_b1_S4406 = 4406;
  localparam test_b1_S4407 = 4407;
  localparam test_b1_S4408 = 4408;
  localparam test_b1_S4409 = 4409;
  localparam test_b1_S4410 = 4410;
  localparam test_b1_S4411 = 4411;
  localparam test_b1_S4412 = 4412;
  localparam test_b1_S4413 = 4413;
  localparam test_b1_S4414 = 4414;
  localparam test_b1_S4415 = 4415;
  localparam test_b1_S4416 = 4416;
  localparam test_b1_S4417 = 4417;
  localparam test_b1_S4418 = 4418;
  localparam test_b1_S4419 = 4419;
  localparam test_b1_S4420 = 4420;
  localparam test_b1_S4421 = 4421;
  localparam test_b1_S4422 = 4422;
  localparam test_b1_S4423 = 4423;
  localparam test_b1_S4424 = 4424;
  localparam test_b1_S4425 = 4425;
  localparam test_b1_S4426 = 4426;
  localparam test_b1_S4427 = 4427;
  localparam test_b1_S4428 = 4428;
  localparam test_b1_S4429 = 4429;
  localparam test_b1_S4430 = 4430;
  localparam test_b1_S4431 = 4431;
  localparam test_b1_S4432 = 4432;
  localparam test_b1_S4433 = 4433;
  localparam test_b1_S4434 = 4434;
  localparam test_b1_S4435 = 4435;
  localparam test_b1_S4436 = 4436;
  localparam test_b1_S4437 = 4437;
  localparam test_b1_S4438 = 4438;
  localparam test_b1_S4439 = 4439;
  localparam test_b1_S4440 = 4440;
  localparam test_b1_S4441 = 4441;
  localparam test_b1_S4442 = 4442;
  localparam test_b1_S4443 = 4443;
  localparam test_b1_S4444 = 4444;
  localparam test_b1_S4445 = 4445;
  localparam test_b1_S4446 = 4446;
  localparam test_b1_S4447 = 4447;
  localparam test_b1_S4448 = 4448;
  localparam test_b1_S4449 = 4449;
  localparam test_b1_S4450 = 4450;
  localparam test_b1_S4451 = 4451;
  localparam test_b1_S4452 = 4452;
  localparam test_b1_S4453 = 4453;
  localparam test_b1_S4454 = 4454;
  localparam test_b1_S4455 = 4455;
  localparam test_b1_S4456 = 4456;
  localparam test_b1_S4457 = 4457;
  localparam test_b1_S4458 = 4458;
  localparam test_b1_S4459 = 4459;
  localparam test_b1_S4460 = 4460;
  localparam test_b1_S4461 = 4461;
  localparam test_b1_S4462 = 4462;
  localparam test_b1_S4463 = 4463;
  localparam test_b1_S4464 = 4464;
  localparam test_b1_S4465 = 4465;
  localparam test_b1_S4466 = 4466;
  localparam test_b1_S4467 = 4467;
  localparam test_b1_S4468 = 4468;
  localparam test_b1_S4469 = 4469;
  localparam test_b1_S4470 = 4470;
  localparam test_b1_S4471 = 4471;
  localparam test_b1_S4472 = 4472;
  localparam test_b1_S4473 = 4473;
  localparam test_b1_S4474 = 4474;
  localparam test_b1_S4475 = 4475;
  localparam test_b1_S4476 = 4476;
  localparam test_b1_S4477 = 4477;
  localparam test_b1_S4478 = 4478;
  localparam test_b1_S4479 = 4479;
  localparam test_b1_S4480 = 4480;
  localparam test_b1_S4481 = 4481;
  localparam test_b1_S4482 = 4482;
  localparam test_b1_S4483 = 4483;
  localparam test_b1_S4484 = 4484;
  localparam test_b1_S4485 = 4485;
  localparam test_b1_S4486 = 4486;
  localparam test_b1_S4487 = 4487;
  localparam test_b1_S4488 = 4488;
  localparam test_b1_S4489 = 4489;
  localparam test_b1_S4490 = 4490;
  localparam test_b1_S4491 = 4491;
  localparam test_b1_S4492 = 4492;
  localparam test_b1_S4493 = 4493;
  localparam test_b1_S4494 = 4494;
  localparam test_b1_S4495 = 4495;
  localparam test_b1_S4496 = 4496;
  localparam test_b1_S4497 = 4497;
  localparam test_b1_S4498 = 4498;
  localparam test_b1_S4499 = 4499;
  localparam test_b1_S4500 = 4500;
  localparam test_b1_S4501 = 4501;
  localparam test_b1_S4502 = 4502;
  localparam test_b1_S4503 = 4503;
  localparam test_b1_S4504 = 4504;
  localparam test_b1_S4505 = 4505;
  localparam test_b1_S4506 = 4506;
  localparam test_b1_S4507 = 4507;
  localparam test_b1_S4508 = 4508;
  localparam test_b1_S4509 = 4509;
  localparam test_b1_S4510 = 4510;
  localparam test_b1_S4511 = 4511;
  localparam test_b1_S4512 = 4512;
  localparam test_b1_S4513 = 4513;
  localparam test_b1_S4514 = 4514;
  localparam test_b1_S4515 = 4515;
  localparam test_b1_S4516 = 4516;
  localparam test_b1_S4517 = 4517;
  localparam test_b1_S4518 = 4518;
  localparam test_b1_S4519 = 4519;
  localparam test_b1_S4520 = 4520;
  localparam test_b1_S4521 = 4521;
  localparam test_b1_S4522 = 4522;
  localparam test_b1_S4523 = 4523;
  localparam test_b1_S4524 = 4524;
  localparam test_b1_S4525 = 4525;
  localparam test_b1_S4526 = 4526;
  localparam test_b1_S4527 = 4527;
  localparam test_b1_S4528 = 4528;
  localparam test_b1_S4529 = 4529;
  localparam test_b1_S4530 = 4530;
  localparam test_b1_S4531 = 4531;
  localparam test_b1_S4532 = 4532;
  localparam test_b1_S4533 = 4533;
  localparam test_b1_S4534 = 4534;
  localparam test_b1_S4535 = 4535;
  localparam test_b1_S4536 = 4536;
  localparam test_b1_S4537 = 4537;
  localparam test_b1_S4538 = 4538;
  localparam test_b1_S4539 = 4539;
  localparam test_b1_S4540 = 4540;
  localparam test_b1_S4541 = 4541;
  localparam test_b1_S4542 = 4542;
  localparam test_b1_S4543 = 4543;
  localparam test_b1_S4544 = 4544;
  localparam test_b1_S4545 = 4545;
  localparam test_b1_S4546 = 4546;
  localparam test_b1_S4547 = 4547;
  localparam test_b1_S4548 = 4548;
  localparam test_b1_S4549 = 4549;
  localparam test_b1_S4550 = 4550;
  localparam test_b1_S4551 = 4551;
  localparam test_b1_S4552 = 4552;
  localparam test_b1_S4553 = 4553;
  localparam test_b1_S4554 = 4554;
  localparam test_b1_S4555 = 4555;
  localparam test_b1_S4556 = 4556;
  localparam test_b1_S4557 = 4557;
  localparam test_b1_S4558 = 4558;
  localparam test_b1_S4559 = 4559;
  localparam test_b1_S4560 = 4560;
  localparam test_b1_S4561 = 4561;
  localparam test_b1_S4562 = 4562;
  localparam test_b1_S4563 = 4563;
  localparam test_b1_S4564 = 4564;
  localparam test_b1_S4565 = 4565;
  localparam test_b1_S4566 = 4566;
  localparam test_b1_S4567 = 4567;
  localparam test_b1_S4568 = 4568;
  localparam test_b1_S4569 = 4569;
  localparam test_b1_S4570 = 4570;
  localparam test_b1_S4571 = 4571;
  localparam test_b1_S4572 = 4572;
  localparam test_b1_S4573 = 4573;
  localparam test_b1_S4574 = 4574;
  localparam test_b1_S4575 = 4575;
  localparam test_b1_S4576 = 4576;
  localparam test_b1_S4577 = 4577;
  localparam test_b1_S4578 = 4578;
  localparam test_b1_S4579 = 4579;
  localparam test_b1_S4580 = 4580;
  localparam test_b1_S4581 = 4581;
  localparam test_b1_S4582 = 4582;
  localparam test_b1_S4583 = 4583;
  localparam test_b1_S4584 = 4584;
  localparam test_b1_S4585 = 4585;
  localparam test_b1_S4586 = 4586;
  localparam test_b1_S4587 = 4587;
  localparam test_b1_S4588 = 4588;
  localparam test_b1_S4589 = 4589;
  localparam test_b1_S4590 = 4590;
  localparam test_b1_S4591 = 4591;
  localparam test_b1_S4592 = 4592;
  localparam test_b1_S4593 = 4593;
  localparam test_b1_S4594 = 4594;
  localparam test_b1_S4595 = 4595;
  localparam test_b1_S4596 = 4596;
  localparam test_b1_S4597 = 4597;
  localparam test_b1_S4598 = 4598;
  localparam test_b1_S4599 = 4599;
  localparam test_b1_S4600 = 4600;
  localparam test_b1_S4601 = 4601;
  localparam test_b1_S4602 = 4602;
  localparam test_b1_S4603 = 4603;
  localparam test_b1_S4604 = 4604;
  localparam test_b1_S4605 = 4605;
  localparam test_b1_S4606 = 4606;
  localparam test_b1_S4607 = 4607;
  localparam test_b1_S4608 = 4608;
  localparam test_b1_S4609 = 4609;
  localparam test_b1_S4610 = 4610;
  localparam test_b1_S4611 = 4611;
  localparam test_b1_S4612 = 4612;
  localparam test_b1_S4613 = 4613;
  localparam test_b1_S4614 = 4614;
  localparam test_b1_S4615 = 4615;
  localparam test_b1_S4616 = 4616;
  localparam test_b1_S4617 = 4617;
  localparam test_b1_S4618 = 4618;
  localparam test_b1_S4619 = 4619;
  localparam test_b1_S4620 = 4620;
  localparam test_b1_S4621 = 4621;
  localparam test_b1_S4622 = 4622;
  localparam test_b1_S4623 = 4623;
  localparam test_b1_S4624 = 4624;
  localparam test_b1_S4625 = 4625;
  localparam test_b1_S4626 = 4626;
  localparam test_b1_S4627 = 4627;
  localparam test_b1_S4628 = 4628;
  localparam test_b1_S4629 = 4629;
  localparam test_b1_S4630 = 4630;
  localparam test_b1_S4631 = 4631;
  localparam test_b1_S4632 = 4632;
  localparam test_b1_S4633 = 4633;
  localparam test_b1_S4634 = 4634;
  localparam test_b1_S4635 = 4635;
  localparam test_b1_S4636 = 4636;
  localparam test_b1_S4637 = 4637;
  localparam test_b1_S4638 = 4638;
  localparam test_b1_S4639 = 4639;
  localparam test_b1_S4640 = 4640;
  localparam test_b1_S4641 = 4641;
  localparam test_b1_S4642 = 4642;
  localparam test_b1_S4643 = 4643;
  localparam test_b1_S4644 = 4644;
  localparam test_b1_S4645 = 4645;
  localparam test_b1_S4646 = 4646;
  localparam test_b1_S4647 = 4647;
  localparam test_b1_S4648 = 4648;
  localparam test_b1_S4649 = 4649;
  localparam test_b1_S4650 = 4650;
  localparam test_b1_S4651 = 4651;
  localparam test_b1_S4652 = 4652;
  localparam test_b1_S4653 = 4653;
  localparam test_b1_S4654 = 4654;
  localparam test_b1_S4655 = 4655;
  localparam test_b1_S4656 = 4656;
  localparam test_b1_S4657 = 4657;
  localparam test_b1_S4658 = 4658;
  localparam test_b1_S4659 = 4659;
  localparam test_b1_S4660 = 4660;
  localparam test_b1_S4661 = 4661;
  localparam test_b1_S4662 = 4662;
  localparam test_b1_S4663 = 4663;
  localparam test_b1_S4664 = 4664;
  localparam test_b1_S4665 = 4665;
  localparam test_b1_S4666 = 4666;
  localparam test_b1_S4667 = 4667;
  localparam test_b1_S4668 = 4668;
  localparam test_b1_S4669 = 4669;
  localparam test_b1_S4670 = 4670;
  localparam test_b1_S4671 = 4671;
  localparam test_b1_S4672 = 4672;
  localparam test_b1_S4673 = 4673;
  localparam test_b1_S4674 = 4674;
  localparam test_b1_S4675 = 4675;
  localparam test_b1_S4676 = 4676;
  localparam test_b1_S4677 = 4677;
  localparam test_b1_S4678 = 4678;
  localparam test_b1_S4679 = 4679;
  localparam test_b1_S4680 = 4680;
  localparam test_b1_S4681 = 4681;
  localparam test_b1_S4682 = 4682;
  localparam test_b1_S4683 = 4683;
  localparam test_b1_S4684 = 4684;
  localparam test_b1_S4685 = 4685;
  localparam test_b1_S4686 = 4686;
  localparam test_b1_S4687 = 4687;
  localparam test_b1_S4688 = 4688;
  localparam test_b1_S4689 = 4689;
  localparam test_b1_S4690 = 4690;
  localparam test_b1_S4691 = 4691;
  localparam test_b1_S4692 = 4692;
  localparam test_b1_S4693 = 4693;
  localparam test_b1_S4694 = 4694;
  localparam test_b1_S4695 = 4695;
  localparam test_b1_S4696 = 4696;
  localparam test_b1_S4697 = 4697;
  localparam test_b1_S4698 = 4698;
  localparam test_b1_S4699 = 4699;
  localparam test_b1_S4700 = 4700;
  localparam test_b1_S4701 = 4701;
  localparam test_b1_S4702 = 4702;
  localparam test_b1_S4703 = 4703;
  localparam test_b1_S4704 = 4704;
  localparam test_b1_S4705 = 4705;
  localparam test_b1_S4706 = 4706;
  localparam test_b1_S4707 = 4707;
  localparam test_b1_S4708 = 4708;
  localparam test_b1_S4709 = 4709;
  localparam test_b1_S4710 = 4710;
  localparam test_b1_S4711 = 4711;
  localparam test_b1_S4712 = 4712;
  localparam test_b1_S4713 = 4713;
  localparam test_b1_S4714 = 4714;
  localparam test_b1_S4715 = 4715;
  localparam test_b1_S4716 = 4716;
  localparam test_b1_S4717 = 4717;
  localparam test_b1_S4718 = 4718;
  localparam test_b1_S4719 = 4719;
  localparam test_b1_S4720 = 4720;
  localparam test_b1_S4721 = 4721;
  localparam test_b1_S4722 = 4722;
  localparam test_b1_S4723 = 4723;
  localparam test_b1_S4724 = 4724;
  localparam test_b1_S4725 = 4725;
  localparam test_b1_S4726 = 4726;
  localparam test_b1_S4727 = 4727;
  localparam test_b1_S4728 = 4728;
  localparam test_b1_S4729 = 4729;
  localparam test_b1_S4730 = 4730;
  localparam test_b1_S4731 = 4731;
  localparam test_b1_S4732 = 4732;
  localparam test_b1_S4733 = 4733;
  localparam test_b1_S4734 = 4734;
  localparam test_b1_S4735 = 4735;
  localparam test_b1_S4736 = 4736;
  localparam test_b1_S4737 = 4737;
  localparam test_b1_S4738 = 4738;
  localparam test_b1_S4739 = 4739;
  localparam test_b1_S4740 = 4740;
  localparam test_b1_S4741 = 4741;
  localparam test_b1_S4742 = 4742;
  localparam test_b1_S4743 = 4743;
  localparam test_b1_S4744 = 4744;
  localparam test_b1_S4745 = 4745;
  localparam test_b1_S4746 = 4746;
  localparam test_b1_S4747 = 4747;
  localparam test_b1_S4748 = 4748;
  localparam test_b1_S4749 = 4749;
  localparam test_b1_S4750 = 4750;
  localparam test_b1_S4751 = 4751;
  localparam test_b1_S4752 = 4752;
  localparam test_b1_S4753 = 4753;
  localparam test_b1_S4754 = 4754;
  localparam test_b1_S4755 = 4755;
  localparam test_b1_S4756 = 4756;
  localparam test_b1_S4757 = 4757;
  localparam test_b1_S4758 = 4758;
  localparam test_b1_S4759 = 4759;
  localparam test_b1_S4760 = 4760;
  localparam test_b1_S4761 = 4761;
  localparam test_b1_S4762 = 4762;
  localparam test_b1_S4763 = 4763;
  localparam test_b1_S4764 = 4764;
  localparam test_b1_S4765 = 4765;
  localparam test_b1_S4766 = 4766;
  localparam test_b1_S4767 = 4767;
  localparam test_b1_S4768 = 4768;
  localparam test_b1_S4769 = 4769;
  localparam test_b1_S4770 = 4770;
  localparam test_b1_S4771 = 4771;
  localparam test_b1_S4772 = 4772;
  localparam test_b1_S4773 = 4773;
  localparam test_b1_S4774 = 4774;
  localparam test_b1_S4775 = 4775;
  localparam test_b1_S4776 = 4776;
  localparam test_b1_S4777 = 4777;
  localparam test_b1_S4778 = 4778;
  localparam test_b1_S4779 = 4779;
  localparam test_b1_S4780 = 4780;
  localparam test_b1_S4781 = 4781;
  localparam test_b1_S4782 = 4782;
  localparam test_b1_S4783 = 4783;
  localparam test_b1_S4784 = 4784;
  localparam test_b1_S4785 = 4785;
  localparam test_b1_S4786 = 4786;
  localparam test_b1_S4787 = 4787;
  localparam test_b1_S4788 = 4788;
  localparam test_b1_S4789 = 4789;
  localparam test_b1_S4790 = 4790;
  localparam test_b1_S4791 = 4791;
  localparam test_b1_S4792 = 4792;
  localparam test_b1_S4793 = 4793;
  localparam test_b1_S4794 = 4794;
  localparam test_b1_S4795 = 4795;
  localparam test_b1_S4796 = 4796;
  localparam test_b1_S4797 = 4797;
  localparam test_b1_S4798 = 4798;
  localparam test_b1_S4799 = 4799;
  localparam test_b1_S4800 = 4800;
  localparam test_b1_S4801 = 4801;
  localparam test_b1_S4802 = 4802;
  localparam test_b1_S4803 = 4803;
  localparam test_b1_S4804 = 4804;
  localparam test_b1_S4805 = 4805;
  localparam test_b1_S4806 = 4806;
  localparam test_b1_S4807 = 4807;
  localparam test_b1_S4808 = 4808;
  localparam test_b1_S4809 = 4809;
  localparam test_b1_S4810 = 4810;
  localparam test_b1_S4811 = 4811;
  localparam test_b1_S4812 = 4812;
  localparam test_b1_S4813 = 4813;
  localparam test_b1_S4814 = 4814;
  localparam test_b1_S4815 = 4815;
  localparam test_b1_S4816 = 4816;
  localparam test_b1_S4817 = 4817;
  localparam test_b1_S4818 = 4818;
  localparam test_b1_S4819 = 4819;
  localparam test_b1_S4820 = 4820;
  localparam test_b1_S4821 = 4821;
  localparam test_b1_S4822 = 4822;
  localparam test_b1_S4823 = 4823;
  localparam test_b1_S4824 = 4824;
  localparam test_b1_S4825 = 4825;
  localparam test_b1_S4826 = 4826;
  localparam test_b1_S4827 = 4827;
  localparam test_b1_S4828 = 4828;
  localparam test_b1_S4829 = 4829;
  localparam test_b1_S4830 = 4830;
  localparam test_b1_S4831 = 4831;
  localparam test_b1_S4832 = 4832;
  localparam test_b1_S4833 = 4833;
  localparam test_b1_S4834 = 4834;
  localparam test_b1_S4835 = 4835;
  localparam test_b1_S4836 = 4836;
  localparam test_b1_S4837 = 4837;
  localparam test_b1_S4838 = 4838;
  localparam test_b1_S4839 = 4839;
  localparam test_b1_S4840 = 4840;
  localparam test_b1_S4841 = 4841;
  localparam test_b1_S4842 = 4842;
  localparam test_b1_S4843 = 4843;
  localparam test_b1_S4844 = 4844;
  localparam test_b1_S4845 = 4845;
  localparam test_b1_S4846 = 4846;
  localparam test_b1_S4847 = 4847;
  localparam test_b1_S4848 = 4848;
  localparam test_b1_S4849 = 4849;
  localparam test_b1_S4850 = 4850;
  localparam test_b1_S4851 = 4851;
  localparam test_b1_S4852 = 4852;
  localparam test_b1_S4853 = 4853;
  localparam test_b1_S4854 = 4854;
  localparam test_b1_S4855 = 4855;
  localparam test_b1_S4856 = 4856;
  localparam test_b1_S4857 = 4857;
  localparam test_b1_S4858 = 4858;
  localparam test_b1_S4859 = 4859;
  localparam test_b1_S4860 = 4860;
  localparam test_b1_S4861 = 4861;
  localparam test_b1_S4862 = 4862;
  localparam test_b1_S4863 = 4863;
  localparam test_b1_S4864 = 4864;
  localparam test_b1_S4865 = 4865;
  localparam test_b1_S4866 = 4866;
  localparam test_b1_S4867 = 4867;
  localparam test_b1_S4868 = 4868;
  localparam test_b1_S4869 = 4869;
  localparam test_b1_S4870 = 4870;
  localparam test_b1_S4871 = 4871;
  localparam test_b1_S4872 = 4872;
  localparam test_b1_S4873 = 4873;
  localparam test_b1_S4874 = 4874;
  localparam test_b1_S4875 = 4875;
  localparam test_b1_S4876 = 4876;
  localparam test_b1_S4877 = 4877;
  localparam test_b1_S4878 = 4878;
  localparam test_b1_S4879 = 4879;
  localparam test_b1_S4880 = 4880;
  localparam test_b1_S4881 = 4881;
  localparam test_b1_S4882 = 4882;
  localparam test_b1_S4883 = 4883;
  localparam test_b1_S4884 = 4884;
  localparam test_b1_S4885 = 4885;
  localparam test_b1_S4886 = 4886;
  localparam test_b1_S4887 = 4887;
  localparam test_b1_S4888 = 4888;
  localparam test_b1_S4889 = 4889;
  localparam test_b1_S4890 = 4890;
  localparam test_b1_S4891 = 4891;
  localparam test_b1_S4892 = 4892;
  localparam test_b1_S4893 = 4893;
  localparam test_b1_S4894 = 4894;
  localparam test_b1_S4895 = 4895;
  localparam test_b1_S4896 = 4896;
  localparam test_b1_S4897 = 4897;
  localparam test_b1_S4898 = 4898;
  localparam test_b1_S4899 = 4899;
  localparam test_b1_S4900 = 4900;
  localparam test_b1_S4901 = 4901;
  localparam test_b1_S4902 = 4902;
  localparam test_b1_S4903 = 4903;
  localparam test_b1_S4904 = 4904;
  localparam test_b1_S4905 = 4905;
  localparam test_b1_S4906 = 4906;
  localparam test_b1_S4907 = 4907;
  localparam test_b1_S4908 = 4908;
  localparam test_b1_S4909 = 4909;
  localparam test_b1_S4910 = 4910;
  localparam test_b1_S4911 = 4911;
  localparam test_b1_S4912 = 4912;
  localparam test_b1_S4913 = 4913;
  localparam test_b1_S4914 = 4914;
  localparam test_b1_S4915 = 4915;
  localparam test_b1_S4916 = 4916;
  localparam test_b1_S4917 = 4917;
  localparam test_b1_S4918 = 4918;
  localparam test_b1_S4919 = 4919;
  localparam test_b1_S4920 = 4920;
  localparam test_b1_S4921 = 4921;
  localparam test_b1_S4922 = 4922;
  localparam test_b1_S4923 = 4923;
  localparam test_b1_S4924 = 4924;
  localparam test_b1_S4925 = 4925;
  localparam test_b1_S4926 = 4926;
  localparam test_b1_S4927 = 4927;
  localparam test_b1_S4928 = 4928;
  localparam test_b1_S4929 = 4929;
  localparam test_b1_S4930 = 4930;
  localparam test_b1_S4931 = 4931;
  localparam test_b1_S4932 = 4932;
  localparam test_b1_S4933 = 4933;
  localparam test_b1_S4934 = 4934;
  localparam test_b1_S4935 = 4935;
  localparam test_b1_S4936 = 4936;
  localparam test_b1_S4937 = 4937;
  localparam test_b1_S4938 = 4938;
  localparam test_b1_S4939 = 4939;
  localparam test_b1_S4940 = 4940;
  localparam test_b1_S4941 = 4941;
  localparam test_b1_S4942 = 4942;
  localparam test_b1_S4943 = 4943;
  localparam test_b1_S4944 = 4944;
  localparam test_b1_S4945 = 4945;
  localparam test_b1_S4946 = 4946;
  localparam test_b1_S4947 = 4947;
  localparam test_b1_S4948 = 4948;
  localparam test_b1_S4949 = 4949;
  localparam test_b1_S4950 = 4950;
  localparam test_b1_S4951 = 4951;
  localparam test_b1_S4952 = 4952;
  localparam test_b1_S4953 = 4953;
  localparam test_b1_S4954 = 4954;
  localparam test_b1_S4955 = 4955;
  localparam test_b1_S4956 = 4956;
  localparam test_b1_S4957 = 4957;
  localparam test_b1_S4958 = 4958;
  localparam test_b1_S4959 = 4959;
  localparam test_b1_S4960 = 4960;
  localparam test_b1_S4961 = 4961;
  localparam test_b1_S4962 = 4962;
  localparam test_b1_S4963 = 4963;
  localparam test_b1_S4964 = 4964;
  localparam test_b1_S4965 = 4965;
  localparam test_b1_S4966 = 4966;
  localparam test_b1_S4967 = 4967;
  localparam test_b1_S4968 = 4968;
  localparam test_b1_S4969 = 4969;
  localparam test_b1_S4970 = 4970;
  localparam test_b1_S4971 = 4971;
  localparam test_b1_S4972 = 4972;
  localparam test_b1_S4973 = 4973;
  localparam test_b1_S4974 = 4974;
  localparam test_b1_S4975 = 4975;
  localparam test_b1_S4976 = 4976;
  localparam test_b1_S4977 = 4977;
  localparam test_b1_S4978 = 4978;
  localparam test_b1_S4979 = 4979;
  localparam test_b1_S4980 = 4980;
  localparam test_b1_S4981 = 4981;
  localparam test_b1_S4982 = 4982;
  localparam test_b1_S4983 = 4983;
  localparam test_b1_S4984 = 4984;
  localparam test_b1_S4985 = 4985;
  localparam test_b1_S4986 = 4986;
  localparam test_b1_S4987 = 4987;
  localparam test_b1_S4988 = 4988;
  localparam test_b1_S4989 = 4989;
  localparam test_b1_S4990 = 4990;
  localparam test_b1_S4991 = 4991;
  localparam test_b1_S4992 = 4992;
  localparam test_b1_S4993 = 4993;
  localparam test_b1_S4994 = 4994;
  localparam test_b1_S4995 = 4995;
  localparam test_b1_S4996 = 4996;
  localparam test_b1_S4997 = 4997;
  localparam test_b1_S4998 = 4998;
  localparam test_b1_S4999 = 4999;
  localparam test_b1_S5000 = 5000;
  localparam test_b1_S5001 = 5001;
  localparam test_b1_S5002 = 5002;
  localparam test_b1_S5003 = 5003;
  localparam test_b1_S5004 = 5004;
  localparam test_b1_S5005 = 5005;
  localparam test_b1_S5006 = 5006;
  localparam test_b1_S5007 = 5007;
  localparam test_b1_S5008 = 5008;
  localparam test_b1_S5009 = 5009;
  localparam test_b1_S5010 = 5010;
  localparam test_b1_S5011 = 5011;
  localparam test_b1_S5012 = 5012;
  localparam test_b1_S5013 = 5013;
  localparam test_b1_S5014 = 5014;
  localparam test_b1_S5015 = 5015;
  localparam test_b1_S5016 = 5016;
  localparam test_b1_S5017 = 5017;
  localparam test_b1_S5018 = 5018;
  localparam test_b1_S5019 = 5019;
  localparam test_b1_S5020 = 5020;
  localparam test_b1_S5021 = 5021;
  localparam test_b1_S5022 = 5022;
  localparam test_b1_S5023 = 5023;
  localparam test_b1_S5024 = 5024;
  localparam test_b1_S5025 = 5025;
  localparam test_b1_S5026 = 5026;
  localparam test_b1_S5027 = 5027;
  localparam test_b1_S5028 = 5028;
  localparam test_b1_S5029 = 5029;
  localparam test_b1_S5030 = 5030;
  localparam test_b1_S5031 = 5031;
  localparam test_b1_S5032 = 5032;
  localparam test_b1_S5033 = 5033;
  localparam test_b1_S5034 = 5034;
  localparam test_b1_S5035 = 5035;
  localparam test_b1_S5036 = 5036;
  localparam test_b1_S5037 = 5037;
  localparam test_b1_S5038 = 5038;
  localparam test_b1_S5039 = 5039;
  localparam test_b1_S5040 = 5040;
  localparam test_b1_S5041 = 5041;
  localparam test_b1_S5042 = 5042;
  localparam test_b1_S5043 = 5043;
  localparam test_b1_S5044 = 5044;
  localparam test_b1_S5045 = 5045;
  localparam test_b1_S5046 = 5046;
  localparam test_b1_S5047 = 5047;
  localparam test_b1_S5048 = 5048;
  localparam test_b1_S5049 = 5049;
  localparam test_b1_S5050 = 5050;
  localparam test_b1_S5051 = 5051;
  localparam test_b1_S5052 = 5052;
  localparam test_b1_S5053 = 5053;
  localparam test_b1_S5054 = 5054;
  localparam test_b1_S5055 = 5055;
  localparam test_b1_S5056 = 5056;
  localparam test_b1_S5057 = 5057;
  localparam test_b1_S5058 = 5058;
  localparam test_b1_S5059 = 5059;
  localparam test_b1_S5060 = 5060;
  localparam test_b1_S5061 = 5061;
  localparam test_b1_S5062 = 5062;
  localparam test_b1_S5063 = 5063;
  localparam test_b1_S5064 = 5064;
  localparam test_b1_S5065 = 5065;
  localparam test_b1_S5066 = 5066;
  localparam test_b1_S5067 = 5067;
  localparam test_b1_S5068 = 5068;
  localparam test_b1_S5069 = 5069;
  localparam test_b1_S5070 = 5070;
  localparam test_b1_S5071 = 5071;
  localparam test_b1_S5072 = 5072;
  localparam test_b1_S5073 = 5073;
  localparam test_b1_S5074 = 5074;
  localparam test_b1_S5075 = 5075;
  localparam test_b1_S5076 = 5076;
  localparam test_b1_S5077 = 5077;
  localparam test_b1_S5078 = 5078;
  localparam test_b1_S5079 = 5079;
  localparam test_b1_S5080 = 5080;
  localparam test_b1_S5081 = 5081;
  localparam test_b1_S5082 = 5082;
  localparam test_b1_S5083 = 5083;
  localparam test_b1_S5084 = 5084;
  localparam test_b1_S5085 = 5085;
  localparam test_b1_S5086 = 5086;
  localparam test_b1_S5087 = 5087;
  localparam test_b1_S5088 = 5088;
  localparam test_b1_S5089 = 5089;
  localparam test_b1_S5090 = 5090;
  localparam test_b1_S5091 = 5091;
  localparam test_b1_S5092 = 5092;
  localparam test_b1_S5093 = 5093;
  localparam test_b1_S5094 = 5094;
  localparam test_b1_S5095 = 5095;
  localparam test_b1_S5096 = 5096;
  localparam test_b1_S5097 = 5097;
  localparam test_b1_S5098 = 5098;
  localparam test_b1_S5099 = 5099;
  localparam test_b1_S5100 = 5100;
  localparam test_b1_S5101 = 5101;
  localparam test_b1_S5102 = 5102;
  localparam test_b1_S5103 = 5103;
  localparam test_b1_S5104 = 5104;
  localparam test_b1_S5105 = 5105;
  localparam test_b1_S5106 = 5106;
  localparam test_b1_S5107 = 5107;
  localparam test_b1_S5108 = 5108;
  localparam test_b1_S5109 = 5109;
  localparam test_b1_S5110 = 5110;
  localparam test_b1_S5111 = 5111;
  localparam test_b1_S5112 = 5112;
  localparam test_b1_S5113 = 5113;
  localparam test_b1_S5114 = 5114;
  localparam test_b1_S5115 = 5115;
  localparam test_b1_S5116 = 5116;
  localparam test_b1_S5117 = 5117;
  localparam test_b1_S5118 = 5118;
  localparam test_b1_S5119 = 5119;
  localparam test_b1_S5120 = 5120;
  localparam test_b1_S5121 = 5121;
  localparam test_b1_S5122 = 5122;
  localparam test_b1_S5123 = 5123;
  localparam test_b1_S5124 = 5124;
  localparam test_b1_S5125 = 5125;
  localparam test_b1_S5126 = 5126;
  localparam test_b1_S5127 = 5127;
  localparam test_b1_S5128 = 5128;
  localparam test_b1_S5129 = 5129;
  localparam test_b1_S5130 = 5130;
  localparam test_b1_S5131 = 5131;
  localparam test_b1_S5132 = 5132;
  localparam test_b1_S5133 = 5133;
  localparam test_b1_S5134 = 5134;
  localparam test_b1_S5135 = 5135;
  localparam test_b1_S5136 = 5136;
  localparam test_b1_S5137 = 5137;
  localparam test_b1_S5138 = 5138;
  localparam test_b1_S5139 = 5139;
  localparam test_b1_S5140 = 5140;
  localparam test_b1_S5141 = 5141;
  localparam test_b1_S5142 = 5142;
  localparam test_b1_S5143 = 5143;
  localparam test_b1_S5144 = 5144;
  localparam test_b1_S5145 = 5145;
  localparam test_b1_S5146 = 5146;
  localparam test_b1_S5147 = 5147;
  localparam test_b1_S5148 = 5148;
  localparam test_b1_S5149 = 5149;
  localparam test_b1_S5150 = 5150;
  localparam test_b1_S5151 = 5151;
  localparam test_b1_S5152 = 5152;
  localparam test_b1_S5153 = 5153;
  localparam test_b1_S5154 = 5154;
  localparam test_b1_S5155 = 5155;
  localparam test_b1_S5156 = 5156;
  localparam test_b1_S5157 = 5157;
  localparam test_b1_S5158 = 5158;
  localparam test_b1_S5159 = 5159;
  localparam test_b1_S5160 = 5160;
  localparam test_b1_S5161 = 5161;
  localparam test_b1_S5162 = 5162;
  localparam test_b1_S5163 = 5163;
  localparam test_b1_S5164 = 5164;
  localparam test_b1_S5165 = 5165;
  localparam test_b1_S5166 = 5166;
  localparam test_b1_S5167 = 5167;
  localparam test_b1_S5168 = 5168;
  localparam test_b1_S5169 = 5169;
  localparam test_b1_S5170 = 5170;
  localparam test_b1_S5171 = 5171;
  localparam test_b1_S5172 = 5172;
  localparam test_b1_S5173 = 5173;
  localparam test_b1_S5174 = 5174;
  localparam test_b1_S5175 = 5175;
  localparam test_b1_S5176 = 5176;
  localparam test_b1_S5177 = 5177;
  localparam test_b1_S5178 = 5178;
  localparam test_b1_S5179 = 5179;
  localparam test_b1_S5180 = 5180;
  localparam test_b1_S5181 = 5181;
  localparam test_b1_S5182 = 5182;
  localparam test_b1_S5183 = 5183;
  localparam test_b1_S5184 = 5184;
  localparam test_b1_S5185 = 5185;
  localparam test_b1_S5186 = 5186;
  localparam test_b1_S5187 = 5187;
  localparam test_b1_S5188 = 5188;
  localparam test_b1_S5189 = 5189;
  localparam test_b1_S5190 = 5190;
  localparam test_b1_S5191 = 5191;
  localparam test_b1_S5192 = 5192;
  localparam test_b1_S5193 = 5193;
  localparam test_b1_S5194 = 5194;
  localparam test_b1_S5195 = 5195;
  localparam test_b1_S5196 = 5196;
  localparam test_b1_S5197 = 5197;
  localparam test_b1_S5198 = 5198;
  localparam test_b1_S5199 = 5199;
  localparam test_b1_S5200 = 5200;
  localparam test_b1_S5201 = 5201;
  localparam test_b1_S5202 = 5202;
  localparam test_b1_S5203 = 5203;
  localparam test_b1_S5204 = 5204;
  localparam test_b1_S5205 = 5205;
  localparam test_b1_S5206 = 5206;
  localparam test_b1_S5207 = 5207;
  localparam test_b1_S5208 = 5208;
  localparam test_b1_S5209 = 5209;
  localparam test_b1_S5210 = 5210;
  localparam test_b1_S5211 = 5211;
  localparam test_b1_S5212 = 5212;
  localparam test_b1_S5213 = 5213;
  localparam test_b1_S5214 = 5214;
  localparam test_b1_S5215 = 5215;
  localparam test_b1_S5216 = 5216;
  localparam test_b1_S5217 = 5217;
  localparam test_b1_S5218 = 5218;
  localparam test_b1_S5219 = 5219;
  localparam test_b1_S5220 = 5220;
  localparam test_b1_S5221 = 5221;
  localparam test_b1_S5222 = 5222;
  localparam test_b1_S5223 = 5223;
  localparam test_b1_S5224 = 5224;
  localparam test_b1_S5225 = 5225;
  localparam test_b1_S5226 = 5226;
  localparam test_b1_S5227 = 5227;
  localparam test_b1_S5228 = 5228;
  localparam test_b1_S5229 = 5229;
  localparam test_b1_S5230 = 5230;
  localparam test_b1_S5231 = 5231;
  localparam test_b1_S5232 = 5232;
  localparam test_b1_S5233 = 5233;
  localparam test_b1_S5234 = 5234;
  localparam test_b1_S5235 = 5235;
  localparam test_b1_S5236 = 5236;
  localparam test_b1_S5237 = 5237;
  localparam test_b1_S5238 = 5238;
  localparam test_b1_S5239 = 5239;
  localparam test_b1_S5240 = 5240;
  localparam test_b1_S5241 = 5241;
  localparam test_b1_S5242 = 5242;
  localparam test_b1_S5243 = 5243;
  localparam test_b1_S5244 = 5244;
  localparam test_b1_S5245 = 5245;
  localparam test_b1_S5246 = 5246;
  localparam test_b1_S5247 = 5247;
  localparam test_b1_S5248 = 5248;
  localparam test_b1_S5249 = 5249;
  localparam test_b1_S5250 = 5250;
  localparam test_b1_S5251 = 5251;
  localparam test_b1_S5252 = 5252;
  localparam test_b1_S5253 = 5253;
  localparam test_b1_S5254 = 5254;
  localparam test_b1_S5255 = 5255;
  localparam test_b1_S5256 = 5256;
  localparam test_b1_S5257 = 5257;
  localparam test_b1_S5258 = 5258;
  localparam test_b1_S5259 = 5259;
  localparam test_b1_S5260 = 5260;
  localparam test_b1_S5261 = 5261;
  localparam test_b1_S5262 = 5262;
  localparam test_b1_S5263 = 5263;
  localparam test_b1_S5264 = 5264;
  localparam test_b1_S5265 = 5265;
  localparam test_b1_S5266 = 5266;
  localparam test_b1_S5267 = 5267;
  localparam test_b1_S5268 = 5268;
  localparam test_b1_S5269 = 5269;
  localparam test_b1_S5270 = 5270;
  localparam test_b1_S5271 = 5271;
  localparam test_b1_S5272 = 5272;
  localparam test_b1_S5273 = 5273;
  localparam test_b1_S5274 = 5274;
  localparam test_b1_S5275 = 5275;
  localparam test_b1_S5276 = 5276;
  localparam test_b1_S5277 = 5277;
  localparam test_b1_S5278 = 5278;
  localparam test_b1_S5279 = 5279;
  localparam test_b1_S5280 = 5280;
  localparam test_b1_S5281 = 5281;
  localparam test_b1_S5282 = 5282;
  localparam test_b1_S5283 = 5283;
  localparam test_b1_S5284 = 5284;
  localparam test_b1_S5285 = 5285;
  localparam test_b1_S5286 = 5286;
  localparam test_b1_S5287 = 5287;
  localparam test_b1_S5288 = 5288;
  localparam test_b1_S5289 = 5289;
  localparam test_b1_S5290 = 5290;
  localparam test_b1_S5291 = 5291;
  localparam test_b1_S5292 = 5292;
  localparam test_b1_S5293 = 5293;
  localparam test_b1_S5294 = 5294;
  localparam test_b1_S5295 = 5295;
  localparam test_b1_S5296 = 5296;
  localparam test_b1_S5297 = 5297;
  localparam test_b1_S5298 = 5298;
  localparam test_b1_S5299 = 5299;
  localparam test_b1_S5300 = 5300;
  localparam test_b1_S5301 = 5301;
  localparam test_b1_S5302 = 5302;
  localparam test_b1_S5303 = 5303;
  localparam test_b1_S5304 = 5304;
  localparam test_b1_S5305 = 5305;
  localparam test_b1_S5306 = 5306;
  localparam test_b1_S5307 = 5307;
  localparam test_b1_S5308 = 5308;
  localparam test_b1_S5309 = 5309;
  localparam test_b1_S5310 = 5310;
  localparam test_b1_S5311 = 5311;
  localparam test_b1_S5312 = 5312;
  localparam test_b1_S5313 = 5313;
  localparam test_b1_S5314 = 5314;
  localparam test_b1_S5315 = 5315;
  localparam test_b1_S5316 = 5316;
  localparam test_b1_S5317 = 5317;
  localparam test_b1_S5318 = 5318;
  localparam test_b1_S5319 = 5319;
  localparam test_b1_S5320 = 5320;
  localparam test_b1_S5321 = 5321;
  localparam test_b1_S5322 = 5322;
  localparam test_b1_S5323 = 5323;
  localparam test_b1_S5324 = 5324;
  localparam test_b1_S5325 = 5325;
  localparam test_b1_S5326 = 5326;
  localparam test_b1_S5327 = 5327;
  localparam test_b1_S5328 = 5328;
  localparam test_b1_S5329 = 5329;
  localparam test_b1_S5330 = 5330;
  localparam test_b1_S5331 = 5331;
  localparam test_b1_S5332 = 5332;
  localparam test_b1_S5333 = 5333;
  localparam test_b1_S5334 = 5334;
  localparam test_b1_S5335 = 5335;
  localparam test_b1_S5336 = 5336;
  localparam test_b1_S5337 = 5337;
  localparam test_b1_S5338 = 5338;
  localparam test_b1_S5339 = 5339;
  localparam test_b1_S5340 = 5340;
  localparam test_b1_S5341 = 5341;
  localparam test_b1_S5342 = 5342;
  localparam test_b1_S5343 = 5343;
  localparam test_b1_S5344 = 5344;
  localparam test_b1_S5345 = 5345;
  localparam test_b1_S5346 = 5346;
  localparam test_b1_S5347 = 5347;
  localparam test_b1_S5348 = 5348;
  localparam test_b1_S5349 = 5349;
  localparam test_b1_S5350 = 5350;
  localparam test_b1_S5351 = 5351;
  localparam test_b1_S5352 = 5352;
  localparam test_b1_S5353 = 5353;
  localparam test_b1_S5354 = 5354;
  localparam test_b1_S5355 = 5355;
  localparam test_b1_S5356 = 5356;
  localparam test_b1_S5357 = 5357;
  localparam test_b1_S5358 = 5358;
  localparam test_b1_S5359 = 5359;
  localparam test_b1_S5360 = 5360;
  localparam test_b1_S5361 = 5361;
  localparam test_b1_S5362 = 5362;
  localparam test_b1_S5363 = 5363;
  localparam test_b1_S5364 = 5364;
  localparam test_b1_S5365 = 5365;
  localparam test_b1_S5366 = 5366;
  localparam test_b1_S5367 = 5367;
  localparam test_b1_S5368 = 5368;
  localparam test_b1_S5369 = 5369;
  localparam test_b1_S5370 = 5370;
  localparam test_b1_S5371 = 5371;
  localparam test_b1_S5372 = 5372;
  localparam test_b1_S5373 = 5373;
  localparam test_b1_S5374 = 5374;
  localparam test_b1_S5375 = 5375;
  localparam test_b1_S5376 = 5376;
  localparam test_b1_S5377 = 5377;
  localparam test_b1_S5378 = 5378;
  localparam test_b1_S5379 = 5379;
  localparam test_b1_S5380 = 5380;
  localparam test_b1_S5381 = 5381;
  localparam test_b1_S5382 = 5382;
  localparam test_b1_S5383 = 5383;
  localparam test_b1_S5384 = 5384;
  localparam test_b1_S5385 = 5385;
  localparam test_b1_S5386 = 5386;
  localparam test_b1_S5387 = 5387;
  localparam test_b1_S5388 = 5388;
  localparam test_b1_S5389 = 5389;
  localparam test_b1_S5390 = 5390;
  localparam test_b1_S5391 = 5391;
  localparam test_b1_S5392 = 5392;
  localparam test_b1_S5393 = 5393;
  localparam test_b1_S5394 = 5394;
  localparam test_b1_S5395 = 5395;
  localparam test_b1_S5396 = 5396;
  localparam test_b1_S5397 = 5397;
  localparam test_b1_S5398 = 5398;
  localparam test_b1_S5399 = 5399;
  localparam test_b1_S5400 = 5400;
  localparam test_b1_S5401 = 5401;
  localparam test_b1_S5402 = 5402;
  localparam test_b1_S5403 = 5403;
  localparam test_b1_S5404 = 5404;
  localparam test_b1_S5405 = 5405;
  localparam test_b1_S5406 = 5406;
  localparam test_b1_S5407 = 5407;
  localparam test_b1_S5408 = 5408;
  localparam test_b1_S5409 = 5409;
  localparam test_b1_S5410 = 5410;
  localparam test_b1_S5411 = 5411;
  localparam test_b1_S5412 = 5412;
  localparam test_b1_S5413 = 5413;
  localparam test_b1_S5414 = 5414;
  localparam test_b1_S5415 = 5415;
  localparam test_b1_S5416 = 5416;
  localparam test_b1_S5417 = 5417;
  localparam test_b1_S5418 = 5418;
  localparam test_b1_S5419 = 5419;
  localparam test_b1_S5420 = 5420;
  localparam test_b1_S5421 = 5421;
  localparam test_b1_S5422 = 5422;
  localparam test_b1_S5423 = 5423;
  localparam test_b1_S5424 = 5424;
  localparam test_b1_S5425 = 5425;
  localparam test_b1_S5426 = 5426;
  localparam test_b1_S5427 = 5427;
  localparam test_b1_S5428 = 5428;
  localparam test_b1_S5429 = 5429;
  localparam test_b1_S5430 = 5430;
  localparam test_b1_S5431 = 5431;
  localparam test_b1_S5432 = 5432;
  localparam test_b1_S5433 = 5433;
  localparam test_b1_S5434 = 5434;
  localparam test_b1_S5435 = 5435;
  localparam test_b1_S5436 = 5436;
  localparam test_b1_S5437 = 5437;
  localparam test_b1_S5438 = 5438;
  localparam test_b1_S5439 = 5439;
  localparam test_b1_S5440 = 5440;
  localparam test_b1_S5441 = 5441;
  localparam test_b1_S5442 = 5442;
  localparam test_b1_S5443 = 5443;
  localparam test_b1_S5444 = 5444;
  localparam test_b1_S5445 = 5445;
  localparam test_b1_S5446 = 5446;
  localparam test_b1_S5447 = 5447;
  localparam test_b1_S5448 = 5448;
  localparam test_b1_S5449 = 5449;
  localparam test_b1_S5450 = 5450;
  localparam test_b1_S5451 = 5451;
  localparam test_b1_S5452 = 5452;
  localparam test_b1_S5453 = 5453;
  localparam test_b1_S5454 = 5454;
  localparam test_b1_S5455 = 5455;
  localparam test_b1_S5456 = 5456;
  localparam test_b1_S5457 = 5457;
  localparam test_b1_S5458 = 5458;
  localparam test_b1_S5459 = 5459;
  localparam test_b1_S5460 = 5460;
  localparam test_b1_S5461 = 5461;
  localparam test_b1_S5462 = 5462;
  localparam test_b1_S5463 = 5463;
  localparam test_b1_S5464 = 5464;
  localparam test_b1_S5465 = 5465;
  localparam test_b1_S5466 = 5466;
  localparam test_b1_S5467 = 5467;
  localparam test_b1_S5468 = 5468;
  localparam test_b1_S5469 = 5469;
  localparam test_b1_S5470 = 5470;
  localparam test_b1_S5471 = 5471;
  localparam test_b1_S5472 = 5472;
  localparam test_b1_S5473 = 5473;
  localparam test_b1_S5474 = 5474;
  localparam test_b1_S5475 = 5475;
  localparam test_b1_S5476 = 5476;
  localparam test_b1_S5477 = 5477;
  localparam test_b1_S5478 = 5478;
  localparam test_b1_S5479 = 5479;
  localparam test_b1_S5480 = 5480;
  localparam test_b1_S5481 = 5481;
  localparam test_b1_S5482 = 5482;
  localparam test_b1_S5483 = 5483;
  localparam test_b1_S5484 = 5484;
  localparam test_b1_S5485 = 5485;
  localparam test_b1_S5486 = 5486;
  localparam test_b1_S5487 = 5487;
  localparam test_b1_S5488 = 5488;
  localparam test_b1_S5489 = 5489;
  localparam test_b1_S5490 = 5490;
  localparam test_b1_S5491 = 5491;
  localparam test_b1_S5492 = 5492;
  localparam test_b1_S5493 = 5493;
  localparam test_b1_S5494 = 5494;
  localparam test_b1_S5495 = 5495;
  localparam test_b1_S5496 = 5496;
  localparam test_b1_S5497 = 5497;
  localparam test_b1_S5498 = 5498;
  localparam test_b1_S5499 = 5499;
  localparam test_b1_S5500 = 5500;
  localparam test_b1_S5501 = 5501;
  localparam test_b1_S5502 = 5502;
  localparam test_b1_S5503 = 5503;
  localparam test_b1_S5504 = 5504;
  localparam test_b1_S5505 = 5505;
  localparam test_b1_S5506 = 5506;
  localparam test_b1_S5507 = 5507;
  localparam test_b1_S5508 = 5508;
  localparam test_b1_S5509 = 5509;
  localparam test_b1_S5510 = 5510;
  localparam test_b1_S5511 = 5511;
  localparam test_b1_S5512 = 5512;
  localparam test_b1_S5513 = 5513;
  localparam test_b1_S5514 = 5514;
  localparam test_b1_S5515 = 5515;
  localparam test_b1_S5516 = 5516;
  localparam test_b1_S5517 = 5517;
  localparam test_b1_S5518 = 5518;
  localparam test_b1_S5519 = 5519;
  localparam test_b1_S5520 = 5520;
  localparam test_b1_S5521 = 5521;
  localparam test_b1_S5522 = 5522;
  localparam test_b1_S5523 = 5523;
  localparam test_b1_S5524 = 5524;
  localparam test_b1_S5525 = 5525;
  localparam test_b1_S5526 = 5526;
  localparam test_b1_S5527 = 5527;
  localparam test_b1_S5528 = 5528;
  localparam test_b1_S5529 = 5529;
  localparam test_b1_S5530 = 5530;
  localparam test_b1_S5531 = 5531;
  localparam test_b1_S5532 = 5532;
  localparam test_b1_S5533 = 5533;
  localparam test_b1_S5534 = 5534;
  localparam test_b1_S5535 = 5535;
  localparam test_b1_S5536 = 5536;
  localparam test_b1_S5537 = 5537;
  localparam test_b1_S5538 = 5538;
  localparam test_b1_S5539 = 5539;
  localparam test_b1_S5540 = 5540;
  localparam test_b1_S5541 = 5541;
  localparam test_b1_S5542 = 5542;
  localparam test_b1_S5543 = 5543;
  localparam test_b1_S5544 = 5544;
  localparam test_b1_S5545 = 5545;
  localparam test_b1_S5546 = 5546;
  localparam test_b1_S5547 = 5547;
  localparam test_b1_S5548 = 5548;
  localparam test_b1_S5549 = 5549;
  localparam test_b1_S5550 = 5550;
  localparam test_b1_S5551 = 5551;
  localparam test_b1_S5552 = 5552;
  localparam test_b1_S5553 = 5553;
  localparam test_b1_S5554 = 5554;
  localparam test_b1_S5555 = 5555;
  localparam test_b1_S5556 = 5556;
  localparam test_b1_S5557 = 5557;
  localparam test_b1_S5558 = 5558;
  localparam test_b1_S5559 = 5559;
  localparam test_b1_S5560 = 5560;
  localparam test_b1_S5561 = 5561;
  localparam test_b1_S5562 = 5562;
  localparam test_b1_S5563 = 5563;
  localparam test_b1_S5564 = 5564;
  localparam test_b1_S5565 = 5565;
  localparam test_b1_S5566 = 5566;
  localparam test_b1_S5567 = 5567;
  localparam test_b1_S5568 = 5568;
  localparam test_b1_S5569 = 5569;
  localparam test_b1_S5570 = 5570;
  localparam test_b1_S5571 = 5571;
  localparam test_b1_S5572 = 5572;
  localparam test_b1_S5573 = 5573;
  localparam test_b1_S5574 = 5574;
  localparam test_b1_S5575 = 5575;
  localparam test_b1_S5576 = 5576;
  localparam test_b1_S5577 = 5577;
  localparam test_b1_S5578 = 5578;
  localparam test_b1_S5579 = 5579;
  localparam test_b1_S5580 = 5580;
  localparam test_b1_S5581 = 5581;
  localparam test_b1_S5582 = 5582;
  localparam test_b1_S5583 = 5583;
  localparam test_b1_S5584 = 5584;
  localparam test_b1_S5585 = 5585;
  localparam test_b1_S5586 = 5586;
  localparam test_b1_S5587 = 5587;
  localparam test_b1_S5588 = 5588;
  localparam test_b1_S5589 = 5589;
  localparam test_b1_S5590 = 5590;
  localparam test_b1_S5591 = 5591;
  localparam test_b1_S5592 = 5592;
  localparam test_b1_S5593 = 5593;
  localparam test_b1_S5594 = 5594;
  localparam test_b1_S5595 = 5595;
  localparam test_b1_S5596 = 5596;
  localparam test_b1_S5597 = 5597;
  localparam test_b1_S5598 = 5598;
  localparam test_b1_S5599 = 5599;
  localparam test_b1_S5600 = 5600;
  localparam test_b1_S5601 = 5601;
  localparam test_b1_S5602 = 5602;
  localparam test_b1_S5603 = 5603;
  localparam test_b1_S5604 = 5604;
  localparam test_b1_S5605 = 5605;
  localparam test_b1_S5606 = 5606;
  localparam test_b1_S5607 = 5607;
  localparam test_b1_S5608 = 5608;
  localparam test_b1_S5609 = 5609;
  localparam test_b1_S5610 = 5610;
  localparam test_b1_S5611 = 5611;
  localparam test_b1_S5612 = 5612;
  localparam test_b1_S5613 = 5613;
  localparam test_b1_S5614 = 5614;
  localparam test_b1_S5615 = 5615;
  localparam test_b1_S5616 = 5616;
  localparam test_b1_S5617 = 5617;
  localparam test_b1_S5618 = 5618;
  localparam test_b1_S5619 = 5619;
  localparam test_b1_S5620 = 5620;
  localparam test_b1_S5621 = 5621;
  localparam test_b1_S5622 = 5622;
  localparam test_b1_S5623 = 5623;
  localparam test_b1_S5624 = 5624;
  localparam test_b1_S5625 = 5625;
  localparam test_b1_S5626 = 5626;
  localparam test_b1_S5627 = 5627;
  localparam test_b1_S5628 = 5628;
  localparam test_b1_S5629 = 5629;
  localparam test_b1_S5630 = 5630;
  localparam test_b1_S5631 = 5631;
  localparam test_b1_S5632 = 5632;
  localparam test_b1_S5633 = 5633;
  localparam test_b1_S5634 = 5634;
  localparam test_b1_S5635 = 5635;
  localparam test_b1_S5636 = 5636;
  localparam test_b1_S5637 = 5637;
  localparam test_b1_S5638 = 5638;
  localparam test_b1_S5639 = 5639;
  localparam test_b1_S5640 = 5640;
  localparam test_b1_S5641 = 5641;
  localparam test_b1_S5642 = 5642;
  localparam test_b1_S5643 = 5643;
  localparam test_b1_S5644 = 5644;
  localparam test_b1_S5645 = 5645;
  localparam test_b1_S5646 = 5646;
  localparam test_b1_S5647 = 5647;
  localparam test_b1_S5648 = 5648;
  localparam test_b1_S5649 = 5649;
  localparam test_b1_S5650 = 5650;
  localparam test_b1_S5651 = 5651;
  localparam test_b1_S5652 = 5652;
  localparam test_b1_S5653 = 5653;
  localparam test_b1_S5654 = 5654;
  localparam test_b1_S5655 = 5655;
  localparam test_b1_S5656 = 5656;
  localparam test_b1_S5657 = 5657;
  localparam test_b1_S5658 = 5658;
  localparam test_b1_S5659 = 5659;
  localparam test_b1_S5660 = 5660;
  localparam test_b1_S5661 = 5661;
  localparam test_b1_S5662 = 5662;
  localparam test_b1_S5663 = 5663;
  localparam test_b1_S5664 = 5664;
  localparam test_b1_S5665 = 5665;
  localparam test_b1_S5666 = 5666;
  localparam test_b1_S5667 = 5667;
  localparam test_b1_S5668 = 5668;
  localparam test_b1_S5669 = 5669;
  localparam test_b1_S5670 = 5670;
  localparam test_b1_S5671 = 5671;
  localparam test_b1_S5672 = 5672;
  localparam test_b1_S5673 = 5673;
  localparam test_b1_S5674 = 5674;
  localparam test_b1_S5675 = 5675;
  localparam test_b1_S5676 = 5676;
  localparam test_b1_S5677 = 5677;
  localparam test_b1_S5678 = 5678;
  localparam test_b1_S5679 = 5679;
  localparam test_b1_S5680 = 5680;
  localparam test_b1_S5681 = 5681;
  localparam test_b1_S5682 = 5682;
  localparam test_b1_S5683 = 5683;
  localparam test_b1_S5684 = 5684;
  localparam test_b1_S5685 = 5685;
  localparam test_b1_S5686 = 5686;
  localparam test_b1_S5687 = 5687;
  localparam test_b1_S5688 = 5688;
  localparam test_b1_S5689 = 5689;
  localparam test_b1_S5690 = 5690;
  localparam test_b1_S5691 = 5691;
  localparam test_b1_S5692 = 5692;
  localparam test_b1_S5693 = 5693;
  localparam test_b1_S5694 = 5694;
  localparam test_b1_S5695 = 5695;
  localparam test_b1_S5696 = 5696;
  localparam test_b1_S5697 = 5697;
  localparam test_b1_S5698 = 5698;
  localparam test_b1_S5699 = 5699;
  localparam test_b1_S5700 = 5700;
  localparam test_b1_S5701 = 5701;
  localparam test_b1_S5702 = 5702;
  localparam test_b1_S5703 = 5703;
  localparam test_b1_S5704 = 5704;
  localparam test_b1_S5705 = 5705;
  localparam test_b1_S5706 = 5706;
  localparam test_b1_S5707 = 5707;
  localparam test_b1_S5708 = 5708;
  localparam test_b1_S5709 = 5709;
  localparam test_b1_S5710 = 5710;
  localparam test_b1_S5711 = 5711;
  localparam test_b1_S5712 = 5712;
  localparam test_b1_S5713 = 5713;
  localparam test_b1_S5714 = 5714;
  localparam test_b1_S5715 = 5715;
  localparam test_b1_S5716 = 5716;
  localparam test_b1_S5717 = 5717;
  localparam test_b1_S5718 = 5718;
  localparam test_b1_S5719 = 5719;
  localparam test_b1_S5720 = 5720;
  localparam test_b1_S5721 = 5721;
  localparam test_b1_S5722 = 5722;
  localparam test_b1_S5723 = 5723;
  localparam test_b1_S5724 = 5724;
  localparam test_b1_S5725 = 5725;
  localparam test_b1_S5726 = 5726;
  localparam test_b1_S5727 = 5727;
  localparam test_b1_S5728 = 5728;
  localparam test_b1_S5729 = 5729;
  localparam test_b1_S5730 = 5730;
  localparam test_b1_S5731 = 5731;
  localparam test_b1_S5732 = 5732;
  localparam test_b1_S5733 = 5733;
  localparam test_b1_S5734 = 5734;
  localparam test_b1_S5735 = 5735;
  localparam test_b1_S5736 = 5736;
  localparam test_b1_S5737 = 5737;
  localparam test_b1_S5738 = 5738;
  localparam test_b1_S5739 = 5739;
  localparam test_b1_S5740 = 5740;
  localparam test_b1_S5741 = 5741;
  localparam test_b1_S5742 = 5742;
  localparam test_b1_S5743 = 5743;
  localparam test_b1_S5744 = 5744;
  localparam test_b1_S5745 = 5745;
  localparam test_b1_S5746 = 5746;
  localparam test_b1_S5747 = 5747;
  localparam test_b1_S5748 = 5748;
  localparam test_b1_S5749 = 5749;
  localparam test_b1_S5750 = 5750;
  localparam test_b1_S5751 = 5751;
  localparam test_b1_S5752 = 5752;
  localparam test_b1_S5753 = 5753;
  localparam test_b1_S5754 = 5754;
  localparam test_b1_S5755 = 5755;
  localparam test_b1_S5756 = 5756;
  localparam test_b1_S5757 = 5757;
  localparam test_b1_S5758 = 5758;
  localparam test_b1_S5759 = 5759;
  localparam test_b1_S5760 = 5760;
  localparam test_b1_S5761 = 5761;
  localparam test_b1_S5762 = 5762;
  localparam test_b1_S5763 = 5763;
  localparam test_b1_S5764 = 5764;
  localparam test_b1_S5765 = 5765;
  localparam test_b1_S5766 = 5766;
  localparam test_b1_S5767 = 5767;
  localparam test_b1_S5768 = 5768;
  localparam test_b1_S5769 = 5769;
  localparam test_b1_S5770 = 5770;
  localparam test_b1_S5771 = 5771;
  localparam test_b1_S5772 = 5772;
  localparam test_b1_S5773 = 5773;
  localparam test_b1_S5774 = 5774;
  localparam test_b1_S5775 = 5775;
  localparam test_b1_S5776 = 5776;
  localparam test_b1_S5777 = 5777;
  localparam test_b1_S5778 = 5778;
  localparam test_b1_S5779 = 5779;
  localparam test_b1_S5780 = 5780;
  localparam test_b1_S5781 = 5781;
  localparam test_b1_S5782 = 5782;
  localparam test_b1_S5783 = 5783;
  localparam test_b1_S5784 = 5784;
  localparam test_b1_S5785 = 5785;
  localparam test_b1_S5786 = 5786;
  localparam test_b1_S5787 = 5787;
  localparam test_b1_S5788 = 5788;
  localparam test_b1_S5789 = 5789;
  localparam test_b1_S5790 = 5790;
  localparam test_b1_S5791 = 5791;
  localparam test_b1_S5792 = 5792;
  localparam test_b1_S5793 = 5793;
  localparam test_b1_S5794 = 5794;
  localparam test_b1_S5795 = 5795;
  localparam test_b1_S5796 = 5796;
  localparam test_b1_S5797 = 5797;
  localparam test_b1_S5798 = 5798;
  localparam test_b1_S5799 = 5799;
  localparam test_b1_S5800 = 5800;
  localparam test_b1_S5801 = 5801;
  localparam test_b1_S5802 = 5802;
  localparam test_b1_S5803 = 5803;
  localparam test_b1_S5804 = 5804;
  localparam test_b1_S5805 = 5805;
  localparam test_b1_S5806 = 5806;
  localparam test_b1_S5807 = 5807;
  localparam test_b1_S5808 = 5808;
  localparam test_b1_S5809 = 5809;
  localparam test_b1_S5810 = 5810;
  localparam test_b1_S5811 = 5811;
  localparam test_b1_S5812 = 5812;
  localparam test_b1_S5813 = 5813;
  localparam test_b1_S5814 = 5814;
  localparam test_b1_S5815 = 5815;
  localparam test_b1_S5816 = 5816;
  localparam test_b1_S5817 = 5817;
  localparam test_b1_S5818 = 5818;
  localparam test_b1_S5819 = 5819;
  localparam test_b1_S5820 = 5820;
  localparam test_b1_S5821 = 5821;
  localparam test_b1_S5822 = 5822;
  localparam test_b1_S5823 = 5823;
  localparam test_b1_S5824 = 5824;
  localparam test_b1_S5825 = 5825;
  localparam test_b1_S5826 = 5826;
  localparam test_b1_S5827 = 5827;
  localparam test_b1_S5828 = 5828;
  localparam test_b1_S5829 = 5829;
  localparam test_b1_S5830 = 5830;
  localparam test_b1_S5831 = 5831;
  localparam test_b1_S5832 = 5832;
  localparam test_b1_S5833 = 5833;
  localparam test_b1_S5834 = 5834;
  localparam test_b1_S5835 = 5835;
  localparam test_b1_S5836 = 5836;
  localparam test_b1_S5837 = 5837;
  localparam test_b1_S5838 = 5838;
  localparam test_b1_S5839 = 5839;
  localparam test_b1_S5840 = 5840;
  localparam test_b1_S5841 = 5841;
  localparam test_b1_S5842 = 5842;
  localparam test_b1_S5843 = 5843;
  localparam test_b1_S5844 = 5844;
  localparam test_b1_S5845 = 5845;
  localparam test_b1_S5846 = 5846;
  localparam test_b1_S5847 = 5847;
  localparam test_b1_S5848 = 5848;
  localparam test_b1_S5849 = 5849;
  localparam test_b1_S5850 = 5850;
  localparam test_b1_S5851 = 5851;
  localparam test_b1_S5852 = 5852;
  localparam test_b1_S5853 = 5853;
  localparam test_b1_S5854 = 5854;
  localparam test_b1_S5855 = 5855;
  localparam test_b1_S5856 = 5856;
  localparam test_b1_S5857 = 5857;
  localparam test_b1_S5858 = 5858;
  localparam test_b1_S5859 = 5859;
  localparam test_b1_S5860 = 5860;
  localparam test_b1_S5861 = 5861;
  localparam test_b1_S5862 = 5862;
  localparam test_b1_S5863 = 5863;
  localparam test_b1_S5864 = 5864;
  localparam test_b1_S5865 = 5865;
  localparam test_b1_S5866 = 5866;
  localparam test_b1_S5867 = 5867;
  localparam test_b1_S5868 = 5868;
  localparam test_b1_S5869 = 5869;
  localparam test_b1_S5870 = 5870;
  localparam test_b1_S5871 = 5871;
  localparam test_b1_S5872 = 5872;
  localparam test_b1_S5873 = 5873;
  localparam test_b1_S5874 = 5874;
  localparam test_b1_S5875 = 5875;
  localparam test_b1_S5876 = 5876;
  localparam test_b1_S5877 = 5877;
  localparam test_b1_S5878 = 5878;
  localparam test_b1_S5879 = 5879;
  localparam test_b1_S5880 = 5880;
  localparam test_b1_S5881 = 5881;
  localparam test_b1_S5882 = 5882;
  localparam test_b1_S5883 = 5883;
  localparam test_b1_S5884 = 5884;
  localparam test_b1_S5885 = 5885;
  localparam test_b1_S5886 = 5886;
  localparam test_b1_S5887 = 5887;
  localparam test_b1_S5888 = 5888;
  localparam test_b1_S5889 = 5889;
  localparam test_b1_S5890 = 5890;
  localparam test_b1_S5891 = 5891;
  localparam test_b1_S5892 = 5892;
  localparam test_b1_S5893 = 5893;
  localparam test_b1_S5894 = 5894;
  localparam test_b1_S5895 = 5895;
  localparam test_b1_S5896 = 5896;
  localparam test_b1_S5897 = 5897;
  localparam test_b1_S5898 = 5898;
  localparam test_b1_S5899 = 5899;
  localparam test_b1_S5900 = 5900;
  localparam test_b1_S5901 = 5901;
  localparam test_b1_S5902 = 5902;
  localparam test_b1_S5903 = 5903;
  localparam test_b1_S5904 = 5904;
  localparam test_b1_S5905 = 5905;
  localparam test_b1_S5906 = 5906;
  localparam test_b1_S5907 = 5907;
  localparam test_b1_S5908 = 5908;
  localparam test_b1_S5909 = 5909;
  localparam test_b1_S5910 = 5910;
  localparam test_b1_S5911 = 5911;
  localparam test_b1_S5912 = 5912;
  localparam test_b1_S5913 = 5913;
  localparam test_b1_S5914 = 5914;
  localparam test_b1_S5915 = 5915;
  localparam test_b1_S5916 = 5916;
  localparam test_b1_S5917 = 5917;
  localparam test_b1_S5918 = 5918;
  localparam test_b1_S5919 = 5919;
  localparam test_b1_S5920 = 5920;
  localparam test_b1_S5921 = 5921;
  localparam test_b1_S5922 = 5922;
  localparam test_b1_S5923 = 5923;
  localparam test_b1_S5924 = 5924;
  localparam test_b1_S5925 = 5925;
  localparam test_b1_S5926 = 5926;
  localparam test_b1_S5927 = 5927;
  localparam test_b1_S5928 = 5928;
  localparam test_b1_S5929 = 5929;
  localparam test_b1_S5930 = 5930;
  localparam test_b1_S5931 = 5931;
  localparam test_b1_S5932 = 5932;
  localparam test_b1_S5933 = 5933;
  localparam test_b1_S5934 = 5934;
  localparam test_b1_S5935 = 5935;
  localparam test_b1_S5936 = 5936;
  localparam test_b1_S5937 = 5937;
  localparam test_b1_S5938 = 5938;
  localparam test_b1_S5939 = 5939;
  localparam test_b1_S5940 = 5940;
  localparam test_b1_S5941 = 5941;
  localparam test_b1_S5942 = 5942;
  localparam test_b1_S5943 = 5943;
  localparam test_b1_S5944 = 5944;
  localparam test_b1_S5945 = 5945;
  localparam test_b1_S5946 = 5946;
  localparam test_b1_S5947 = 5947;
  localparam test_b1_S5948 = 5948;
  localparam test_b1_S5949 = 5949;
  localparam test_b1_S5950 = 5950;
  localparam test_b1_S5951 = 5951;
  localparam test_b1_S5952 = 5952;
  localparam test_b1_S5953 = 5953;
  localparam test_b1_S5954 = 5954;
  localparam test_b1_S5955 = 5955;
  localparam test_b1_S5956 = 5956;
  localparam test_b1_S5957 = 5957;
  localparam test_b1_S5958 = 5958;
  localparam test_b1_S5959 = 5959;
  localparam test_b1_S5960 = 5960;
  localparam test_b1_S5961 = 5961;
  localparam test_b1_S5962 = 5962;
  localparam test_b1_S5963 = 5963;
  localparam test_b1_S5964 = 5964;
  localparam test_b1_S5965 = 5965;
  localparam test_b1_S5966 = 5966;
  localparam test_b1_S5967 = 5967;
  localparam test_b1_S5968 = 5968;
  localparam test_b1_S5969 = 5969;
  localparam test_b1_S5970 = 5970;
  localparam test_b1_S5971 = 5971;
  localparam test_b1_S5972 = 5972;
  localparam test_b1_S5973 = 5973;
  localparam test_b1_S5974 = 5974;
  localparam test_b1_S5975 = 5975;
  localparam test_b1_S5976 = 5976;
  localparam test_b1_S5977 = 5977;
  localparam test_b1_S5978 = 5978;
  localparam test_b1_S5979 = 5979;
  localparam test_b1_S5980 = 5980;
  localparam test_b1_S5981 = 5981;
  localparam test_b1_S5982 = 5982;
  localparam test_b1_S5983 = 5983;
  localparam test_b1_S5984 = 5984;
  localparam test_b1_S5985 = 5985;
  localparam test_b1_S5986 = 5986;
  localparam test_b1_S5987 = 5987;
  localparam test_b1_S5988 = 5988;
  localparam test_b1_S5989 = 5989;
  localparam test_b1_S5990 = 5990;
  localparam test_b1_S5991 = 5991;
  localparam test_b1_S5992 = 5992;
  localparam test_b1_S5993 = 5993;
  localparam test_b1_S5994 = 5994;
  localparam test_b1_S5995 = 5995;
  localparam test_b1_S5996 = 5996;
  localparam test_b1_S5997 = 5997;
  localparam test_b1_S5998 = 5998;
  localparam test_b1_S5999 = 5999;
  localparam test_b1_S6000 = 6000;
  localparam test_b1_S6001 = 6001;
  localparam test_b1_S6002 = 6002;
  localparam test_b1_S6003 = 6003;
  localparam test_b1_S6004 = 6004;
  localparam test_b1_S6005 = 6005;
  localparam test_b1_S6006 = 6006;
  localparam test_b1_S6007 = 6007;
  localparam test_b1_S6008 = 6008;
  localparam test_b1_S6009 = 6009;
  localparam test_b1_S6010 = 6010;
  localparam test_b1_S6011 = 6011;
  localparam test_b1_S6012 = 6012;
  localparam test_b1_S6013 = 6013;
  localparam test_b1_S6014 = 6014;
  localparam test_b1_S6015 = 6015;
  localparam test_b1_S6016 = 6016;
  localparam test_b1_S6017 = 6017;
  localparam test_b1_S6018 = 6018;
  localparam test_b1_S6019 = 6019;
  localparam test_b1_S6020 = 6020;
  localparam test_b1_S6021 = 6021;
  localparam test_b1_S6022 = 6022;
  localparam test_b1_S6023 = 6023;
  localparam test_b1_S6024 = 6024;
  localparam test_b1_S6025 = 6025;
  localparam test_b1_S6026 = 6026;
  localparam test_b1_S6027 = 6027;
  localparam test_b1_S6028 = 6028;
  localparam test_b1_S6029 = 6029;
  localparam test_b1_S6030 = 6030;
  localparam test_b1_S6031 = 6031;
  localparam test_b1_S6032 = 6032;
  localparam test_b1_S6033 = 6033;
  localparam test_b1_S6034 = 6034;
  localparam test_b1_S6035 = 6035;
  localparam test_b1_S6036 = 6036;
  localparam test_b1_S6037 = 6037;
  localparam test_b1_S6038 = 6038;
  localparam test_b1_S6039 = 6039;
  localparam test_b1_S6040 = 6040;
  localparam test_b1_S6041 = 6041;
  localparam test_b1_S6042 = 6042;
  localparam test_b1_S6043 = 6043;
  localparam test_b1_S6044 = 6044;
  localparam test_b1_S6045 = 6045;
  localparam test_b1_S6046 = 6046;
  localparam test_b1_S6047 = 6047;
  localparam test_b1_S6048 = 6048;
  localparam test_b1_S6049 = 6049;
  localparam test_b1_S6050 = 6050;
  localparam test_b1_S6051 = 6051;
  localparam test_b1_S6052 = 6052;
  localparam test_b1_S6053 = 6053;
  localparam test_b1_S6054 = 6054;
  localparam test_b1_S6055 = 6055;
  localparam test_b1_S6056 = 6056;
  localparam test_b1_S6057 = 6057;
  localparam test_b1_S6058 = 6058;
  localparam test_b1_S6059 = 6059;
  localparam test_b1_S6060 = 6060;
  localparam test_b1_S6061 = 6061;
  localparam test_b1_S6062 = 6062;
  localparam test_b1_S6063 = 6063;
  localparam test_b1_S6064 = 6064;
  localparam test_b1_S6065 = 6065;
  localparam test_b1_S6066 = 6066;
  localparam test_b1_S6067 = 6067;
  localparam test_b1_S6068 = 6068;
  localparam test_b1_S6069 = 6069;
  localparam test_b1_S6070 = 6070;
  localparam test_b1_S6071 = 6071;
  localparam test_b1_S6072 = 6072;
  localparam test_b1_S6073 = 6073;
  localparam test_b1_S6074 = 6074;
  localparam test_b1_S6075 = 6075;
  localparam test_b1_S6076 = 6076;
  localparam test_b1_S6077 = 6077;
  localparam test_b1_S6078 = 6078;
  localparam test_b1_S6079 = 6079;
  localparam test_b1_S6080 = 6080;
  localparam test_b1_S6081 = 6081;
  localparam test_b1_S6082 = 6082;
  localparam test_b1_S6083 = 6083;
  localparam test_b1_S6084 = 6084;
  localparam test_b1_S6085 = 6085;
  localparam test_b1_S6086 = 6086;
  localparam test_b1_S6087 = 6087;
  localparam test_b1_S6088 = 6088;
  localparam test_b1_S6089 = 6089;
  localparam test_b1_S6090 = 6090;
  localparam test_b1_S6091 = 6091;
  localparam test_b1_S6092 = 6092;
  localparam test_b1_S6093 = 6093;
  localparam test_b1_S6094 = 6094;
  localparam test_b1_S6095 = 6095;
  localparam test_b1_S6096 = 6096;
  localparam test_b1_S6097 = 6097;
  localparam test_b1_S6098 = 6098;
  localparam test_b1_S6099 = 6099;
  localparam test_b1_S6100 = 6100;
  localparam test_b1_S6101 = 6101;
  localparam test_b1_S6102 = 6102;
  localparam test_b1_S6103 = 6103;
  localparam test_b1_S6104 = 6104;
  localparam test_b1_S6105 = 6105;
  localparam test_b1_S6106 = 6106;
  localparam test_b1_S6107 = 6107;
  localparam test_b1_S6108 = 6108;
  localparam test_b1_S6109 = 6109;
  localparam test_b1_S6110 = 6110;
  localparam test_b1_S6111 = 6111;
  localparam test_b1_S6112 = 6112;
  localparam test_b1_S6113 = 6113;
  localparam test_b1_S6114 = 6114;
  localparam test_b1_S6115 = 6115;
  localparam test_b1_S6116 = 6116;
  localparam test_b1_S6117 = 6117;
  localparam test_b1_S6118 = 6118;
  localparam test_b1_S6119 = 6119;
  localparam test_b1_S6120 = 6120;
  localparam test_b1_S6121 = 6121;
  localparam test_b1_S6122 = 6122;
  localparam test_b1_S6123 = 6123;
  localparam test_b1_S6124 = 6124;
  localparam test_b1_S6125 = 6125;
  localparam test_b1_S6126 = 6126;
  localparam test_b1_S6127 = 6127;
  localparam test_b1_S6128 = 6128;
  localparam test_b1_S6129 = 6129;
  localparam test_b1_S6130 = 6130;
  localparam test_b1_S6131 = 6131;
  localparam test_b1_S6132 = 6132;
  localparam test_b1_S6133 = 6133;
  localparam test_b1_S6134 = 6134;
  localparam test_b1_S6135 = 6135;
  localparam test_b1_S6136 = 6136;
  localparam test_b1_S6137 = 6137;
  localparam test_b1_S6138 = 6138;
  localparam test_b1_S6139 = 6139;
  localparam test_b1_S6140 = 6140;
  localparam test_b1_S6141 = 6141;
  localparam test_b1_S6142 = 6142;
  localparam test_b1_S6143 = 6143;
  localparam test_b1_S6144 = 6144;
  localparam test_b1_S6145 = 6145;
  localparam test_b1_S6146 = 6146;
  localparam test_b1_S6147 = 6147;
  localparam test_b1_S6148 = 6148;
  localparam test_b1_S6149 = 6149;
  localparam test_b1_S6150 = 6150;
  localparam test_b1_S6151 = 6151;
  localparam test_b1_S6152 = 6152;
  localparam test_b1_S6153 = 6153;
  localparam test_b1_S6154 = 6154;
  localparam test_b1_S6155 = 6155;
  localparam test_b1_S6156 = 6156;
  localparam test_b1_S6157 = 6157;
  localparam test_b1_S6158 = 6158;
  localparam test_b1_S6159 = 6159;
  localparam test_b1_S6160 = 6160;
  localparam test_b1_S6161 = 6161;
  localparam test_b1_S6162 = 6162;
  localparam test_b1_S6163 = 6163;
  localparam test_b1_S6164 = 6164;
  localparam test_b1_S6165 = 6165;
  localparam test_b1_S6166 = 6166;
  localparam test_b1_S6167 = 6167;
  localparam test_b1_S6168 = 6168;
  localparam test_b1_S6169 = 6169;
  localparam test_b1_S6170 = 6170;
  localparam test_b1_S6171 = 6171;
  localparam test_b1_S6172 = 6172;
  localparam test_b1_S6173 = 6173;
  localparam test_b1_S6174 = 6174;
  localparam test_b1_S6175 = 6175;
  localparam test_b1_S6176 = 6176;
  localparam test_b1_S6177 = 6177;
  localparam test_b1_S6178 = 6178;
  localparam test_b1_S6179 = 6179;
  localparam test_b1_S6180 = 6180;
  localparam test_b1_S6181 = 6181;
  localparam test_b1_S6182 = 6182;
  localparam test_b1_S6183 = 6183;
  localparam test_b1_S6184 = 6184;
  localparam test_b1_S6185 = 6185;
  localparam test_b1_S6186 = 6186;
  localparam test_b1_S6187 = 6187;
  localparam test_b1_S6188 = 6188;
  localparam test_b1_S6189 = 6189;
  localparam test_b1_S6190 = 6190;
  localparam test_b1_S6191 = 6191;
  localparam test_b1_S6192 = 6192;
  localparam test_b1_S6193 = 6193;
  localparam test_b1_S6194 = 6194;
  localparam test_b1_S6195 = 6195;
  localparam test_b1_S6196 = 6196;
  localparam test_b1_S6197 = 6197;
  localparam test_b1_S6198 = 6198;
  localparam test_b1_S6199 = 6199;
  localparam test_b1_S6200 = 6200;
  localparam test_b1_S6201 = 6201;
  localparam test_b1_S6202 = 6202;
  localparam test_b1_S6203 = 6203;
  localparam test_b1_S6204 = 6204;
  localparam test_b1_S6205 = 6205;
  localparam test_b1_S6206 = 6206;
  localparam test_b1_S6207 = 6207;
  localparam test_b1_S6208 = 6208;
  localparam test_b1_S6209 = 6209;
  localparam test_b1_S6210 = 6210;
  localparam test_b1_S6211 = 6211;
  localparam test_b1_S6212 = 6212;
  localparam test_b1_S6213 = 6213;
  localparam test_b1_S6214 = 6214;
  localparam test_b1_S6215 = 6215;
  localparam test_b1_S6216 = 6216;
  localparam test_b1_S6217 = 6217;
  localparam test_b1_S6218 = 6218;
  localparam test_b1_S6219 = 6219;
  localparam test_b1_S6220 = 6220;
  localparam test_b1_S6221 = 6221;
  localparam test_b1_S6222 = 6222;
  localparam test_b1_S6223 = 6223;
  localparam test_b1_S6224 = 6224;
  localparam test_b1_S6225 = 6225;
  localparam test_b1_S6226 = 6226;
  localparam test_b1_S6227 = 6227;
  localparam test_b1_S6228 = 6228;
  localparam test_b1_S6229 = 6229;
  localparam test_b1_S6230 = 6230;
  localparam test_b1_S6231 = 6231;
  localparam test_b1_S6232 = 6232;
  localparam test_b1_S6233 = 6233;
  localparam test_b1_S6234 = 6234;
  localparam test_b1_S6235 = 6235;
  localparam test_b1_S6236 = 6236;
  localparam test_b1_S6237 = 6237;
  localparam test_b1_S6238 = 6238;
  localparam test_b1_S6239 = 6239;
  localparam test_b1_S6240 = 6240;
  localparam test_b1_S6241 = 6241;
  localparam test_b1_S6242 = 6242;
  localparam test_b1_S6243 = 6243;
  localparam test_b1_S6244 = 6244;
  localparam test_b1_S6245 = 6245;
  localparam test_b1_S6246 = 6246;
  localparam test_b1_S6247 = 6247;
  localparam test_b1_S6248 = 6248;
  localparam test_b1_S6249 = 6249;
  localparam test_b1_S6250 = 6250;
  localparam test_b1_S6251 = 6251;
  localparam test_b1_S6252 = 6252;
  localparam test_b1_S6253 = 6253;
  localparam test_b1_S6254 = 6254;
  localparam test_b1_S6255 = 6255;
  localparam test_b1_S6256 = 6256;
  localparam test_b1_S6257 = 6257;
  localparam test_b1_S6258 = 6258;
  localparam test_b1_S6259 = 6259;
  localparam test_b1_S6260 = 6260;
  localparam test_b1_S6261 = 6261;
  localparam test_b1_S6262 = 6262;
  localparam test_b1_S6263 = 6263;
  localparam test_b1_S6264 = 6264;
  localparam test_b1_S6265 = 6265;
  localparam test_b1_S6266 = 6266;
  localparam test_b1_S6267 = 6267;
  localparam test_b1_S6268 = 6268;
  localparam test_b1_S6269 = 6269;
  localparam test_b1_S6270 = 6270;
  localparam test_b1_S6271 = 6271;
  localparam test_b1_S6272 = 6272;
  localparam test_b1_S6273 = 6273;
  localparam test_b1_S6274 = 6274;
  localparam test_b1_S6275 = 6275;
  localparam test_b1_S6276 = 6276;
  localparam test_b1_S6277 = 6277;
  localparam test_b1_S6278 = 6278;
  localparam test_b1_S6279 = 6279;
  localparam test_b1_S6280 = 6280;
  localparam test_b1_S6281 = 6281;
  localparam test_b1_S6282 = 6282;
  localparam test_b1_S6283 = 6283;
  localparam test_b1_S6284 = 6284;
  localparam test_b1_S6285 = 6285;
  localparam test_b1_S6286 = 6286;
  localparam test_b1_S6287 = 6287;
  localparam test_b1_S6288 = 6288;
  localparam test_b1_S6289 = 6289;
  localparam test_b1_S6290 = 6290;
  localparam test_b1_S6291 = 6291;
  localparam test_b1_S6292 = 6292;
  localparam test_b1_S6293 = 6293;
  localparam test_b1_S6294 = 6294;
  localparam test_b1_S6295 = 6295;
  localparam test_b1_S6296 = 6296;
  localparam test_b1_S6297 = 6297;
  localparam test_b1_S6298 = 6298;
  localparam test_b1_S6299 = 6299;
  localparam test_b1_S6300 = 6300;
  localparam test_b1_S6301 = 6301;
  localparam test_b1_S6302 = 6302;
  localparam test_b1_S6303 = 6303;
  localparam test_b1_S6304 = 6304;
  localparam test_b1_S6305 = 6305;
  localparam test_b1_S6306 = 6306;
  localparam test_b1_S6307 = 6307;
  localparam test_b1_S6308 = 6308;
  localparam test_b1_S6309 = 6309;
  localparam test_b1_S6310 = 6310;
  localparam test_b1_S6311 = 6311;
  localparam test_b1_S6312 = 6312;
  localparam test_b1_S6313 = 6313;
  localparam test_b1_S6314 = 6314;
  localparam test_b1_S6315 = 6315;
  localparam test_b1_S6316 = 6316;
  localparam test_b1_S6317 = 6317;
  localparam test_b1_S6318 = 6318;
  localparam test_b1_S6319 = 6319;
  localparam test_b1_S6320 = 6320;
  localparam test_b1_S6321 = 6321;
  localparam test_b1_S6322 = 6322;
  localparam test_b1_S6323 = 6323;
  localparam test_b1_S6324 = 6324;
  localparam test_b1_S6325 = 6325;
  localparam test_b1_S6326 = 6326;
  localparam test_b1_S6327 = 6327;
  localparam test_b1_S6328 = 6328;
  localparam test_b1_S6329 = 6329;
  localparam test_b1_S6330 = 6330;
  localparam test_b1_S6331 = 6331;
  localparam test_b1_S6332 = 6332;
  localparam test_b1_S6333 = 6333;
  localparam test_b1_S6334 = 6334;
  localparam test_b1_S6335 = 6335;
  localparam test_b1_S6336 = 6336;
  localparam test_b1_S6337 = 6337;
  localparam test_b1_S6338 = 6338;
  localparam test_b1_S6339 = 6339;
  localparam test_b1_S6340 = 6340;
  localparam test_b1_S6341 = 6341;
  localparam test_b1_S6342 = 6342;
  localparam test_b1_S6343 = 6343;
  localparam test_b1_S6344 = 6344;
  localparam test_b1_S6345 = 6345;
  localparam test_b1_S6346 = 6346;
  localparam test_b1_S6347 = 6347;
  localparam test_b1_S6348 = 6348;
  localparam test_b1_S6349 = 6349;
  localparam test_b1_S6350 = 6350;
  localparam test_b1_S6351 = 6351;
  localparam test_b1_S6352 = 6352;
  localparam test_b1_S6353 = 6353;
  localparam test_b1_S6354 = 6354;
  localparam test_b1_S6355 = 6355;
  localparam test_b1_S6356 = 6356;
  localparam test_b1_S6357 = 6357;
  localparam test_b1_S6358 = 6358;
  localparam test_b1_S6359 = 6359;
  localparam test_b1_S6360 = 6360;
  localparam test_b1_S6361 = 6361;
  localparam test_b1_S6362 = 6362;
  localparam test_b1_S6363 = 6363;
  localparam test_b1_S6364 = 6364;
  localparam test_b1_S6365 = 6365;
  localparam test_b1_S6366 = 6366;
  localparam test_b1_S6367 = 6367;
  localparam test_b1_S6368 = 6368;
  localparam test_b1_S6369 = 6369;
  localparam test_b1_S6370 = 6370;
  localparam test_b1_S6371 = 6371;
  localparam test_b1_S6372 = 6372;
  localparam test_b1_S6373 = 6373;
  localparam test_b1_S6374 = 6374;
  localparam test_b1_S6375 = 6375;
  localparam test_b1_S6376 = 6376;
  localparam test_b1_S6377 = 6377;
  localparam test_b1_S6378 = 6378;
  localparam test_b1_S6379 = 6379;
  localparam test_b1_S6380 = 6380;
  localparam test_b1_S6381 = 6381;
  localparam test_b1_S6382 = 6382;
  localparam test_b1_S6383 = 6383;
  localparam test_b1_S6384 = 6384;
  localparam test_b1_S6385 = 6385;
  localparam test_b1_S6386 = 6386;
  localparam test_b1_S6387 = 6387;
  localparam test_b1_S6388 = 6388;
  localparam test_b1_S6389 = 6389;
  localparam test_b1_S6390 = 6390;
  localparam test_b1_S6391 = 6391;
  localparam test_b1_S6392 = 6392;
  localparam test_b1_S6393 = 6393;
  localparam test_b1_S6394 = 6394;
  localparam test_b1_S6395 = 6395;
  localparam test_b1_S6396 = 6396;
  localparam test_b1_S6397 = 6397;
  localparam test_b1_S6398 = 6398;
  localparam test_b1_S6399 = 6399;
  localparam test_b1_S6400 = 6400;
  localparam test_b1_S6401 = 6401;
  localparam test_b1_S6402 = 6402;
  localparam test_b1_S6403 = 6403;
  localparam test_b1_S6404 = 6404;
  localparam test_b1_S6405 = 6405;
  localparam test_b1_S6406 = 6406;
  localparam test_b1_S6407 = 6407;
  localparam test_b1_S6408 = 6408;
  localparam test_b1_S6409 = 6409;
  localparam test_b1_S6410 = 6410;
  localparam test_b1_S6411 = 6411;
  localparam test_b1_S6412 = 6412;
  localparam test_b1_S6413 = 6413;
  localparam test_b1_S6414 = 6414;
  localparam test_b1_S6415 = 6415;
  localparam test_b1_S6416 = 6416;
  localparam test_b1_S6417 = 6417;
  localparam test_b1_S6418 = 6418;
  localparam test_b1_S6419 = 6419;
  localparam test_b1_S6420 = 6420;
  localparam test_b1_S6421 = 6421;
  localparam test_b1_S6422 = 6422;
  localparam test_b1_S6423 = 6423;
  localparam test_b1_S6424 = 6424;
  localparam test_b1_S6425 = 6425;
  localparam test_b1_S6426 = 6426;
  localparam test_b1_S6427 = 6427;
  localparam test_b1_S6428 = 6428;
  localparam test_b1_S6429 = 6429;
  localparam test_b1_S6430 = 6430;
  localparam test_b1_S6431 = 6431;
  localparam test_b1_S6432 = 6432;
  localparam test_b1_S6433 = 6433;
  localparam test_b1_S6434 = 6434;
  localparam test_b1_S6435 = 6435;
  localparam test_b1_S6436 = 6436;
  localparam test_b1_S6437 = 6437;
  localparam test_b1_S6438 = 6438;
  localparam test_b1_S6439 = 6439;
  localparam test_b1_S6440 = 6440;
  localparam test_b1_S6441 = 6441;
  localparam test_b1_S6442 = 6442;
  localparam test_b1_S6443 = 6443;
  localparam test_b1_S6444 = 6444;
  localparam test_b1_S6445 = 6445;
  localparam test_b1_S6446 = 6446;
  localparam test_b1_S6447 = 6447;
  localparam test_b1_S6448 = 6448;
  localparam test_b1_S6449 = 6449;
  localparam test_b1_S6450 = 6450;
  localparam test_b1_S6451 = 6451;
  localparam test_b1_S6452 = 6452;
  localparam test_b1_S6453 = 6453;
  localparam test_b1_S6454 = 6454;
  localparam test_b1_S6455 = 6455;
  localparam test_b1_S6456 = 6456;
  localparam test_b1_S6457 = 6457;
  localparam test_b1_S6458 = 6458;
  localparam test_b1_S6459 = 6459;
  localparam test_b1_S6460 = 6460;
  localparam test_b1_S6461 = 6461;
  localparam test_b1_S6462 = 6462;
  localparam test_b1_S6463 = 6463;
  localparam test_b1_S6464 = 6464;
  localparam test_b1_S6465 = 6465;
  localparam test_b1_S6466 = 6466;
  localparam test_b1_S6467 = 6467;
  localparam test_b1_S6468 = 6468;
  localparam test_b1_S6469 = 6469;
  localparam test_b1_S6470 = 6470;
  localparam test_b1_S6471 = 6471;
  localparam test_b1_S6472 = 6472;
  localparam test_b1_S6473 = 6473;
  localparam test_b1_S6474 = 6474;
  localparam test_b1_S6475 = 6475;
  localparam test_b1_S6476 = 6476;
  localparam test_b1_S6477 = 6477;
  localparam test_b1_S6478 = 6478;
  localparam test_b1_S6479 = 6479;
  localparam test_b1_S6480 = 6480;
  localparam test_b1_S6481 = 6481;
  localparam test_b1_S6482 = 6482;
  localparam test_b1_S6483 = 6483;
  localparam test_b1_S6484 = 6484;
  localparam test_b1_S6485 = 6485;
  localparam test_b1_S6486 = 6486;
  localparam test_b1_S6487 = 6487;
  localparam test_b1_S6488 = 6488;
  localparam test_b1_S6489 = 6489;
  localparam test_b1_S6490 = 6490;
  localparam test_b1_S6491 = 6491;
  localparam test_b1_S6492 = 6492;
  localparam test_b1_S6493 = 6493;
  localparam test_b1_S6494 = 6494;
  localparam test_b1_S6495 = 6495;
  localparam test_b1_S6496 = 6496;
  localparam test_b1_S6497 = 6497;
  localparam test_b1_S6498 = 6498;
  localparam test_b1_S6499 = 6499;
  localparam test_b1_S6500 = 6500;
  localparam test_b1_S6501 = 6501;
  localparam test_b1_S6502 = 6502;
  localparam test_b1_S6503 = 6503;
  localparam test_b1_S6504 = 6504;
  localparam test_b1_S6505 = 6505;
  localparam test_b1_S6506 = 6506;
  localparam test_b1_S6507 = 6507;
  localparam test_b1_S6508 = 6508;
  localparam test_b1_S6509 = 6509;
  localparam test_b1_S6510 = 6510;
  localparam test_b1_S6511 = 6511;
  localparam test_b1_S6512 = 6512;
  localparam test_b1_S6513 = 6513;
  localparam test_b1_S6514 = 6514;
  localparam test_b1_S6515 = 6515;
  localparam test_b1_S6516 = 6516;
  localparam test_b1_S6517 = 6517;
  localparam test_b1_S6518 = 6518;
  localparam test_b1_S6519 = 6519;
  localparam test_b1_S6520 = 6520;
  localparam test_b1_S6521 = 6521;
  localparam test_b1_S6522 = 6522;
  localparam test_b1_S6523 = 6523;
  localparam test_b1_S6524 = 6524;
  localparam test_b1_S6525 = 6525;
  localparam test_b1_S6526 = 6526;
  localparam test_b1_S6527 = 6527;
  localparam test_b1_S6528 = 6528;
  localparam test_b1_S6529 = 6529;
  localparam test_b1_S6530 = 6530;
  localparam test_b1_S6531 = 6531;
  localparam test_b1_S6532 = 6532;
  localparam test_b1_S6533 = 6533;
  localparam test_b1_S6534 = 6534;
  localparam test_b1_S6535 = 6535;
  localparam test_b1_S6536 = 6536;
  localparam test_b1_S6537 = 6537;
  localparam test_b1_S6538 = 6538;
  localparam test_b1_S6539 = 6539;
  localparam test_b1_S6540 = 6540;
  localparam test_b1_S6541 = 6541;
  localparam test_b1_S6542 = 6542;
  localparam test_b1_S6543 = 6543;
  localparam test_b1_S6544 = 6544;
  localparam test_b1_S6545 = 6545;
  localparam test_b1_S6546 = 6546;
  localparam test_b1_S6547 = 6547;
  localparam test_b1_S6548 = 6548;
  localparam test_b1_S6549 = 6549;
  localparam test_b1_S6550 = 6550;
  localparam test_b1_S6551 = 6551;
  localparam test_b1_S6552 = 6552;
  localparam test_b1_S6553 = 6553;
  localparam test_b1_S6554 = 6554;
  localparam test_b1_S6555 = 6555;
  localparam test_b1_S6556 = 6556;
  localparam test_b1_S6557 = 6557;
  localparam test_b1_S6558 = 6558;
  localparam test_b1_S6559 = 6559;
  localparam test_b1_S6560 = 6560;
  localparam test_b1_S6561 = 6561;
  localparam test_b1_S6562 = 6562;
  localparam test_b1_S6563 = 6563;
  localparam test_b1_S6564 = 6564;
  localparam test_b1_S6565 = 6565;
  localparam test_b1_S6566 = 6566;
  localparam test_b1_S6567 = 6567;
  localparam test_b1_S6568 = 6568;
  localparam test_b1_S6569 = 6569;
  localparam test_b1_S6570 = 6570;
  localparam test_b1_S6571 = 6571;
  localparam test_b1_S6572 = 6572;
  localparam test_b1_S6573 = 6573;
  localparam test_b1_S6574 = 6574;
  localparam test_b1_S6575 = 6575;
  localparam test_b1_S6576 = 6576;
  localparam test_b1_S6577 = 6577;
  localparam test_b1_S6578 = 6578;
  localparam test_b1_S6579 = 6579;
  localparam test_b1_S6580 = 6580;
  localparam test_b1_S6581 = 6581;
  localparam test_b1_S6582 = 6582;
  localparam test_b1_S6583 = 6583;
  localparam test_b1_S6584 = 6584;
  localparam test_b1_S6585 = 6585;
  localparam test_b1_S6586 = 6586;
  localparam test_b1_S6587 = 6587;
  localparam test_b1_S6588 = 6588;
  localparam test_b1_S6589 = 6589;
  localparam test_b1_S6590 = 6590;
  localparam test_b1_S6591 = 6591;
  localparam test_b1_S6592 = 6592;
  localparam test_b1_S6593 = 6593;
  localparam test_b1_S6594 = 6594;
  localparam test_b1_S6595 = 6595;
  localparam test_b1_S6596 = 6596;
  localparam test_b1_S6597 = 6597;
  localparam test_b1_S6598 = 6598;
  localparam test_b1_S6599 = 6599;
  localparam test_b1_S6600 = 6600;
  localparam test_b1_S6601 = 6601;
  localparam test_b1_S6602 = 6602;
  localparam test_b1_S6603 = 6603;
  localparam test_b1_S6604 = 6604;
  localparam test_b1_S6605 = 6605;
  localparam test_b1_S6606 = 6606;
  localparam test_b1_S6607 = 6607;
  localparam test_b1_S6608 = 6608;
  localparam test_b1_S6609 = 6609;
  localparam test_b1_S6610 = 6610;
  localparam test_b1_S6611 = 6611;
  localparam test_b1_S6612 = 6612;
  localparam test_b1_S6613 = 6613;
  localparam test_b1_S6614 = 6614;
  localparam test_b1_S6615 = 6615;
  localparam test_b1_S6616 = 6616;
  localparam test_b1_S6617 = 6617;
  localparam test_b1_S6618 = 6618;
  localparam test_b1_S6619 = 6619;
  localparam test_b1_S6620 = 6620;
  localparam test_b1_S6621 = 6621;
  localparam test_b1_S6622 = 6622;
  localparam test_b1_S6623 = 6623;
  localparam test_b1_S6624 = 6624;
  localparam test_b1_S6625 = 6625;
  localparam test_b1_S6626 = 6626;
  localparam test_b1_S6627 = 6627;
  localparam test_b1_S6628 = 6628;
  localparam test_b1_S6629 = 6629;
  localparam test_b1_S6630 = 6630;
  localparam test_b1_S6631 = 6631;
  localparam test_b1_S6632 = 6632;
  localparam test_b1_S6633 = 6633;
  localparam test_b1_S6634 = 6634;
  localparam test_b1_S6635 = 6635;
  localparam test_b1_S6636 = 6636;
  localparam test_b1_S6637 = 6637;
  localparam test_b1_S6638 = 6638;
  localparam test_b1_S6639 = 6639;
  localparam test_b1_S6640 = 6640;
  localparam test_b1_S6641 = 6641;
  localparam test_b1_S6642 = 6642;
  localparam test_b1_S6643 = 6643;
  localparam test_b1_S6644 = 6644;
  localparam test_b1_S6645 = 6645;
  localparam test_b1_S6646 = 6646;
  localparam test_b1_S6647 = 6647;
  localparam test_b1_S6648 = 6648;
  localparam test_b1_S6649 = 6649;
  localparam test_b1_S6650 = 6650;
  localparam test_b1_S6651 = 6651;
  localparam test_b1_S6652 = 6652;
  localparam test_b1_S6653 = 6653;
  localparam test_b1_S6654 = 6654;
  localparam test_b1_S6655 = 6655;
  localparam test_b1_S6656 = 6656;
  localparam test_b1_S6657 = 6657;
  localparam test_b1_S6658 = 6658;
  localparam test_b1_S6659 = 6659;
  localparam test_b1_S6660 = 6660;
  localparam test_b1_S6661 = 6661;
  localparam test_b1_S6662 = 6662;
  localparam test_b1_S6663 = 6663;
  localparam test_b1_S6664 = 6664;
  localparam test_b1_S6665 = 6665;
  localparam test_b1_S6666 = 6666;
  localparam test_b1_S6667 = 6667;
  localparam test_b1_S6668 = 6668;
  localparam test_b1_S6669 = 6669;
  localparam test_b1_S6670 = 6670;
  localparam test_b1_S6671 = 6671;
  localparam test_b1_S6672 = 6672;
  localparam test_b1_S6673 = 6673;
  localparam test_b1_S6674 = 6674;
  localparam test_b1_S6675 = 6675;
  localparam test_b1_S6676 = 6676;
  localparam test_b1_S6677 = 6677;
  localparam test_b1_S6678 = 6678;
  localparam test_b1_S6679 = 6679;
  localparam test_b1_S6680 = 6680;
  localparam test_b1_S6681 = 6681;
  localparam test_b1_S6682 = 6682;
  localparam test_b1_S6683 = 6683;
  localparam test_b1_S6684 = 6684;
  localparam test_b1_S6685 = 6685;
  localparam test_b1_S6686 = 6686;
  localparam test_b1_S6687 = 6687;
  localparam test_b1_S6688 = 6688;
  localparam test_b1_S6689 = 6689;
  localparam test_b1_S6690 = 6690;
  localparam test_b1_S6691 = 6691;
  localparam test_b1_S6692 = 6692;
  localparam test_b1_S6693 = 6693;
  localparam test_b1_S6694 = 6694;
  localparam test_b1_S6695 = 6695;
  localparam test_b1_S6696 = 6696;
  localparam test_b1_S6697 = 6697;
  localparam test_b1_S6698 = 6698;
  localparam test_b1_S6699 = 6699;
  localparam test_b1_S6700 = 6700;
  localparam test_b1_S6701 = 6701;
  localparam test_b1_S6702 = 6702;
  localparam test_b1_S6703 = 6703;
  localparam test_b1_S6704 = 6704;
  localparam test_b1_S6705 = 6705;
  localparam test_b1_S6706 = 6706;
  localparam test_b1_S6707 = 6707;
  localparam test_b1_S6708 = 6708;
  localparam test_b1_S6709 = 6709;
  localparam test_b1_S6710 = 6710;
  localparam test_b1_S6711 = 6711;
  localparam test_b1_S6712 = 6712;
  localparam test_b1_S6713 = 6713;
  localparam test_b1_S6714 = 6714;
  localparam test_b1_S6715 = 6715;
  localparam test_b1_S6716 = 6716;
  localparam test_b1_S6717 = 6717;
  localparam test_b1_S6718 = 6718;
  localparam test_b1_S6719 = 6719;
  localparam test_b1_S6720 = 6720;
  localparam test_b1_S6721 = 6721;
  localparam test_b1_S6722 = 6722;
  localparam test_b1_S6723 = 6723;
  localparam test_b1_S6724 = 6724;
  localparam test_b1_S6725 = 6725;
  localparam test_b1_S6726 = 6726;
  localparam test_b1_S6727 = 6727;
  localparam test_b1_S6728 = 6728;
  localparam test_b1_S6729 = 6729;
  localparam test_b1_S6730 = 6730;
  localparam test_b1_S6731 = 6731;
  localparam test_b1_S6732 = 6732;
  localparam test_b1_S6733 = 6733;
  localparam test_b1_S6734 = 6734;
  localparam test_b1_S6735 = 6735;
  localparam test_b1_S6736 = 6736;
  localparam test_b1_S6737 = 6737;
  localparam test_b1_S6738 = 6738;
  localparam test_b1_S6739 = 6739;
  localparam test_b1_S6740 = 6740;
  localparam test_b1_S6741 = 6741;
  localparam test_b1_S6742 = 6742;
  localparam test_b1_S6743 = 6743;
  localparam test_b1_S6744 = 6744;
  localparam test_b1_S6745 = 6745;
  localparam test_b1_S6746 = 6746;
  localparam test_b1_S6747 = 6747;
  localparam test_b1_S6748 = 6748;
  localparam test_b1_S6749 = 6749;
  localparam test_b1_S6750 = 6750;
  localparam test_b1_S6751 = 6751;
  localparam test_b1_S6752 = 6752;
  localparam test_b1_S6753 = 6753;
  localparam test_b1_S6754 = 6754;
  localparam test_b1_S6755 = 6755;
  localparam test_b1_S6756 = 6756;
  localparam test_b1_S6757 = 6757;
  localparam test_b1_S6758 = 6758;
  localparam test_b1_S6759 = 6759;
  localparam test_b1_S6760 = 6760;
  localparam test_b1_S6761 = 6761;
  localparam test_b1_S6762 = 6762;
  localparam test_b1_S6763 = 6763;
  localparam test_b1_S6764 = 6764;
  localparam test_b1_S6765 = 6765;
  localparam test_b1_S6766 = 6766;
  localparam test_b1_S6767 = 6767;
  localparam test_b1_S6768 = 6768;
  localparam test_b1_S6769 = 6769;
  localparam test_b1_S6770 = 6770;
  localparam test_b1_S6771 = 6771;
  localparam test_b1_S6772 = 6772;
  localparam test_b1_S6773 = 6773;
  localparam test_b1_S6774 = 6774;
  localparam test_b1_S6775 = 6775;
  localparam test_b1_S6776 = 6776;
  localparam test_b1_S6777 = 6777;
  localparam test_b1_S6778 = 6778;
  localparam test_b1_S6779 = 6779;
  localparam test_b1_S6780 = 6780;
  localparam test_b1_S6781 = 6781;
  localparam test_b1_S6782 = 6782;
  localparam test_b1_S6783 = 6783;
  localparam test_b1_S6784 = 6784;
  localparam test_b1_S6785 = 6785;
  localparam test_b1_S6786 = 6786;
  localparam test_b1_S6787 = 6787;
  localparam test_b1_S6788 = 6788;
  localparam test_b1_S6789 = 6789;
  localparam test_b1_S6790 = 6790;
  localparam test_b1_S6791 = 6791;
  localparam test_b1_S6792 = 6792;
  localparam test_b1_S6793 = 6793;
  localparam test_b1_S6794 = 6794;
  localparam test_b1_S6795 = 6795;
  localparam test_b1_S6796 = 6796;
  localparam test_b1_S6797 = 6797;
  localparam test_b1_S6798 = 6798;
  localparam test_b1_S6799 = 6799;
  localparam test_b1_S6800 = 6800;
  localparam test_b1_S6801 = 6801;
  localparam test_b1_S6802 = 6802;
  localparam test_b1_S6803 = 6803;
  localparam test_b1_S6804 = 6804;
  localparam test_b1_S6805 = 6805;
  localparam test_b1_S6806 = 6806;
  localparam test_b1_S6807 = 6807;
  localparam test_b1_S6808 = 6808;
  localparam test_b1_S6809 = 6809;
  localparam test_b1_S6810 = 6810;
  localparam test_b1_S6811 = 6811;
  localparam test_b1_S6812 = 6812;
  localparam test_b1_S6813 = 6813;
  localparam test_b1_S6814 = 6814;
  localparam test_b1_S6815 = 6815;
  localparam test_b1_S6816 = 6816;
  localparam test_b1_S6817 = 6817;
  localparam test_b1_S6818 = 6818;
  localparam test_b1_S6819 = 6819;
  localparam test_b1_S6820 = 6820;
  localparam test_b1_S6821 = 6821;
  localparam test_b1_S6822 = 6822;
  localparam test_b1_S6823 = 6823;
  localparam test_b1_S6824 = 6824;
  localparam test_b1_S6825 = 6825;
  localparam test_b1_S6826 = 6826;
  localparam test_b1_S6827 = 6827;
  localparam test_b1_S6828 = 6828;
  localparam test_b1_S6829 = 6829;
  localparam test_b1_S6830 = 6830;
  localparam test_b1_S6831 = 6831;
  localparam test_b1_S6832 = 6832;
  localparam test_b1_S6833 = 6833;
  localparam test_b1_S6834 = 6834;
  localparam test_b1_S6835 = 6835;
  localparam test_b1_S6836 = 6836;
  localparam test_b1_S6837 = 6837;
  localparam test_b1_S6838 = 6838;
  localparam test_b1_S6839 = 6839;
  localparam test_b1_S6840 = 6840;
  localparam test_b1_S6841 = 6841;
  localparam test_b1_S6842 = 6842;
  localparam test_b1_S6843 = 6843;
  localparam test_b1_S6844 = 6844;
  localparam test_b1_S6845 = 6845;
  localparam test_b1_S6846 = 6846;
  localparam test_b1_S6847 = 6847;
  localparam test_b1_S6848 = 6848;
  localparam test_b1_S6849 = 6849;
  localparam test_b1_S6850 = 6850;
  localparam test_b1_S6851 = 6851;
  localparam test_b1_S6852 = 6852;
  localparam test_b1_S6853 = 6853;
  localparam test_b1_S6854 = 6854;
  localparam test_b1_S6855 = 6855;
  localparam test_b1_S6856 = 6856;
  localparam test_b1_S6857 = 6857;
  localparam test_b1_S6858 = 6858;
  localparam test_b1_S6859 = 6859;
  localparam test_b1_S6860 = 6860;
  localparam test_b1_S6861 = 6861;
  localparam test_b1_S6862 = 6862;
  localparam test_b1_S6863 = 6863;
  localparam test_b1_S6864 = 6864;
  localparam test_b1_S6865 = 6865;
  localparam test_b1_S6866 = 6866;
  localparam test_b1_S6867 = 6867;
  localparam test_b1_S6868 = 6868;
  localparam test_b1_S6869 = 6869;
  localparam test_b1_S6870 = 6870;
  localparam test_b1_S6871 = 6871;
  localparam test_b1_S6872 = 6872;
  localparam test_b1_S6873 = 6873;
  localparam test_b1_S6874 = 6874;
  localparam test_b1_S6875 = 6875;
  localparam test_b1_S6876 = 6876;
  localparam test_b1_S6877 = 6877;
  localparam test_b1_S6878 = 6878;
  localparam test_b1_S6879 = 6879;
  localparam test_b1_S6880 = 6880;
  localparam test_b1_S6881 = 6881;
  localparam test_b1_S6882 = 6882;
  localparam test_b1_S6883 = 6883;
  localparam test_b1_S6884 = 6884;
  localparam test_b1_S6885 = 6885;
  localparam test_b1_S6886 = 6886;
  localparam test_b1_S6887 = 6887;
  localparam test_b1_S6888 = 6888;
  localparam test_b1_S6889 = 6889;
  localparam test_b1_S6890 = 6890;
  localparam test_b1_S6891 = 6891;
  localparam test_b1_S6892 = 6892;
  localparam test_b1_S6893 = 6893;
  localparam test_b1_S6894 = 6894;
  localparam test_b1_S6895 = 6895;
  localparam test_b1_S6896 = 6896;
  localparam test_b1_S6897 = 6897;
  localparam test_b1_S6898 = 6898;
  localparam test_b1_S6899 = 6899;
  localparam test_b1_S6900 = 6900;
  localparam test_b1_S6901 = 6901;
  localparam test_b1_S6902 = 6902;
  localparam test_b1_S6903 = 6903;
  localparam test_b1_S6904 = 6904;
  localparam test_b1_S6905 = 6905;
  localparam test_b1_S6906 = 6906;
  localparam test_b1_S6907 = 6907;
  localparam test_b1_S6908 = 6908;
  localparam test_b1_S6909 = 6909;
  localparam test_b1_S6910 = 6910;
  localparam test_b1_S6911 = 6911;
  localparam test_b1_S6912 = 6912;
  localparam test_b1_S6913 = 6913;
  localparam test_b1_S6914 = 6914;
  localparam test_b1_S6915 = 6915;
  localparam test_b1_S6916 = 6916;
  localparam test_b1_S6917 = 6917;
  localparam test_b1_S6918 = 6918;
  localparam test_b1_S6919 = 6919;
  localparam test_b1_S6920 = 6920;
  localparam test_b1_S6921 = 6921;
  localparam test_b1_S6922 = 6922;
  localparam test_b1_S6923 = 6923;
  localparam test_b1_S6924 = 6924;
  localparam test_b1_S6925 = 6925;
  localparam test_b1_S6926 = 6926;
  localparam test_b1_S6927 = 6927;
  localparam test_b1_S6928 = 6928;
  localparam test_b1_S6929 = 6929;
  localparam test_b1_S6930 = 6930;
  localparam test_b1_S6931 = 6931;
  localparam test_b1_S6932 = 6932;
  localparam test_b1_S6933 = 6933;
  localparam test_b1_S6934 = 6934;
  localparam test_b1_S6935 = 6935;
  localparam test_b1_S6936 = 6936;
  localparam test_b1_S6937 = 6937;
  localparam test_b1_S6938 = 6938;
  localparam test_b1_S6939 = 6939;
  localparam test_b1_S6940 = 6940;
  localparam test_b1_S6941 = 6941;
  localparam test_b1_S6942 = 6942;
  localparam test_b1_S6943 = 6943;
  localparam test_b1_S6944 = 6944;
  localparam test_b1_S6945 = 6945;
  localparam test_b1_S6946 = 6946;
  localparam test_b1_S6947 = 6947;
  localparam test_b1_S6948 = 6948;
  localparam test_b1_S6949 = 6949;
  localparam test_b1_S6950 = 6950;
  localparam test_b1_S6951 = 6951;
  localparam test_b1_S6952 = 6952;
  localparam test_b1_S6953 = 6953;
  localparam test_b1_S6954 = 6954;
  localparam test_b1_S6955 = 6955;
  localparam test_b1_S6956 = 6956;
  localparam test_b1_S6957 = 6957;
  localparam test_b1_S6958 = 6958;
  localparam test_b1_S6959 = 6959;
  localparam test_b1_S6960 = 6960;
  localparam test_b1_S6961 = 6961;
  localparam test_b1_S6962 = 6962;
  localparam test_b1_S6963 = 6963;
  localparam test_b1_S6964 = 6964;
  localparam test_b1_S6965 = 6965;
  localparam test_b1_S6966 = 6966;
  localparam test_b1_S6967 = 6967;
  localparam test_b1_S6968 = 6968;
  localparam test_b1_S6969 = 6969;
  localparam test_b1_S6970 = 6970;
  localparam test_b1_S6971 = 6971;
  localparam test_b1_S6972 = 6972;
  localparam test_b1_S6973 = 6973;
  localparam test_b1_S6974 = 6974;
  localparam test_b1_S6975 = 6975;
  localparam test_b1_S6976 = 6976;
  localparam test_b1_S6977 = 6977;
  localparam test_b1_S6978 = 6978;
  localparam test_b1_S6979 = 6979;
  localparam test_b1_S6980 = 6980;
  localparam test_b1_S6981 = 6981;
  localparam test_b1_S6982 = 6982;
  localparam test_b1_S6983 = 6983;
  localparam test_b1_S6984 = 6984;
  localparam test_b1_S6985 = 6985;
  localparam test_b1_S6986 = 6986;
  localparam test_b1_S6987 = 6987;
  localparam test_b1_S6988 = 6988;
  localparam test_b1_S6989 = 6989;
  localparam test_b1_S6990 = 6990;
  localparam test_b1_S6991 = 6991;
  localparam test_b1_S6992 = 6992;
  localparam test_b1_S6993 = 6993;
  localparam test_b1_S6994 = 6994;
  localparam test_b1_S6995 = 6995;
  localparam test_b1_S6996 = 6996;
  localparam test_b1_S6997 = 6997;
  localparam test_b1_S6998 = 6998;
  localparam test_b1_S6999 = 6999;
  localparam test_b1_S7000 = 7000;
  localparam test_b1_S7001 = 7001;
  localparam test_b1_S7002 = 7002;
  localparam test_b1_S7003 = 7003;
  localparam test_b1_S7004 = 7004;
  localparam test_b1_S7005 = 7005;
  localparam test_b1_S7006 = 7006;
  localparam test_b1_S7007 = 7007;
  localparam test_b1_S7008 = 7008;
  localparam test_b1_S7009 = 7009;
  localparam test_b1_S7010 = 7010;
  localparam test_b1_S7011 = 7011;
  localparam test_b1_S7012 = 7012;
  localparam test_b1_S7013 = 7013;
  localparam test_b1_S7014 = 7014;
  localparam test_b1_S7015 = 7015;
  localparam test_b1_S7016 = 7016;
  localparam test_b1_S7017 = 7017;
  localparam test_b1_S7018 = 7018;
  localparam test_b1_S7019 = 7019;
  localparam test_b1_S7020 = 7020;
  localparam test_b1_S7021 = 7021;
  localparam test_b1_S7022 = 7022;
  localparam test_b1_S7023 = 7023;
  localparam test_b1_S7024 = 7024;
  localparam test_b1_S7025 = 7025;
  localparam test_b1_S7026 = 7026;
  localparam test_b1_S7027 = 7027;
  localparam test_b1_S7028 = 7028;
  localparam test_b1_S7029 = 7029;
  localparam test_b1_S7030 = 7030;
  localparam test_b1_S7031 = 7031;
  localparam test_b1_S7032 = 7032;
  localparam test_b1_S7033 = 7033;
  localparam test_b1_S7034 = 7034;
  localparam test_b1_S7035 = 7035;
  localparam test_b1_S7036 = 7036;
  localparam test_b1_S7037 = 7037;
  localparam test_b1_S7038 = 7038;
  localparam test_b1_S7039 = 7039;
  localparam test_b1_S7040 = 7040;
  localparam test_b1_S7041 = 7041;
  localparam test_b1_S7042 = 7042;
  localparam test_b1_S7043 = 7043;
  localparam test_b1_S7044 = 7044;
  localparam test_b1_S7045 = 7045;
  localparam test_b1_S7046 = 7046;
  localparam test_b1_S7047 = 7047;
  localparam test_b1_S7048 = 7048;
  localparam test_b1_S7049 = 7049;
  localparam test_b1_S7050 = 7050;
  localparam test_b1_S7051 = 7051;
  localparam test_b1_S7052 = 7052;
  localparam test_b1_S7053 = 7053;
  localparam test_b1_S7054 = 7054;
  localparam test_b1_S7055 = 7055;
  localparam test_b1_S7056 = 7056;
  localparam test_b1_S7057 = 7057;
  localparam test_b1_S7058 = 7058;
  localparam test_b1_S7059 = 7059;
  localparam test_b1_S7060 = 7060;
  localparam test_b1_S7061 = 7061;
  localparam test_b1_S7062 = 7062;
  localparam test_b1_S7063 = 7063;
  localparam test_b1_S7064 = 7064;
  localparam test_b1_S7065 = 7065;
  localparam test_b1_S7066 = 7066;
  localparam test_b1_S7067 = 7067;
  localparam test_b1_S7068 = 7068;
  localparam test_b1_S7069 = 7069;
  localparam test_b1_S7070 = 7070;
  localparam test_b1_S7071 = 7071;
  localparam test_b1_S7072 = 7072;
  localparam test_b1_S7073 = 7073;
  localparam test_b1_S7074 = 7074;
  localparam test_b1_S7075 = 7075;
  localparam test_b1_S7076 = 7076;
  localparam test_b1_S7077 = 7077;
  localparam test_b1_S7078 = 7078;
  localparam test_b1_S7079 = 7079;
  localparam test_b1_S7080 = 7080;
  localparam test_b1_S7081 = 7081;
  localparam test_b1_S7082 = 7082;
  localparam test_b1_S7083 = 7083;
  localparam test_b1_S7084 = 7084;
  localparam test_b1_S7085 = 7085;
  localparam test_b1_S7086 = 7086;
  localparam test_b1_S7087 = 7087;
  localparam test_b1_S7088 = 7088;
  localparam test_b1_S7089 = 7089;
  localparam test_b1_S7090 = 7090;
  localparam test_b1_S7091 = 7091;
  localparam test_b1_S7092 = 7092;
  localparam test_b1_S7093 = 7093;
  localparam test_b1_S7094 = 7094;
  localparam test_b1_S7095 = 7095;
  localparam test_b1_S7096 = 7096;
  localparam test_b1_S7097 = 7097;
  localparam test_b1_S7098 = 7098;
  localparam test_b1_S7099 = 7099;
  localparam test_b1_S7100 = 7100;
  localparam test_b1_S7101 = 7101;
  localparam test_b1_S7102 = 7102;
  localparam test_b1_S7103 = 7103;
  localparam test_b1_S7104 = 7104;
  localparam test_b1_S7105 = 7105;
  localparam test_b1_S7106 = 7106;
  localparam test_b1_S7107 = 7107;
  localparam test_b1_S7108 = 7108;
  localparam test_b1_S7109 = 7109;
  localparam test_b1_S7110 = 7110;
  localparam test_b1_S7111 = 7111;
  localparam test_b1_S7112 = 7112;
  localparam test_b1_S7113 = 7113;
  localparam test_b1_S7114 = 7114;
  localparam test_b1_S7115 = 7115;
  localparam test_b1_S7116 = 7116;
  localparam test_b1_S7117 = 7117;
  localparam test_b1_S7118 = 7118;
  localparam test_b1_S7119 = 7119;
  localparam test_b1_S7120 = 7120;
  localparam test_b1_S7121 = 7121;
  localparam test_b1_S7122 = 7122;
  localparam test_b1_S7123 = 7123;
  localparam test_b1_S7124 = 7124;
  localparam test_b1_S7125 = 7125;
  localparam test_b1_S7126 = 7126;
  localparam test_b1_S7127 = 7127;
  localparam test_b1_S7128 = 7128;
  localparam test_b1_S7129 = 7129;
  localparam test_b1_S7130 = 7130;
  localparam test_b1_S7131 = 7131;
  localparam test_b1_S7132 = 7132;
  localparam test_b1_S7133 = 7133;
  localparam test_b1_S7134 = 7134;
  localparam test_b1_S7135 = 7135;
  localparam test_b1_S7136 = 7136;
  localparam test_b1_S7137 = 7137;
  localparam test_b1_S7138 = 7138;
  localparam test_b1_S7139 = 7139;
  localparam test_b1_S7140 = 7140;
  localparam test_b1_S7141 = 7141;
  localparam test_b1_S7142 = 7142;
  localparam test_b1_S7143 = 7143;
  localparam test_b1_S7144 = 7144;
  localparam test_b1_S7145 = 7145;
  localparam test_b1_S7146 = 7146;
  localparam test_b1_S7147 = 7147;
  localparam test_b1_S7148 = 7148;
  localparam test_b1_S7149 = 7149;
  localparam test_b1_S7150 = 7150;
  localparam test_b1_S7151 = 7151;
  localparam test_b1_S7152 = 7152;
  localparam test_b1_S7153 = 7153;
  localparam test_b1_S7154 = 7154;
  localparam test_b1_S7155 = 7155;
  localparam test_b1_S7156 = 7156;
  localparam test_b1_S7157 = 7157;
  localparam test_b1_S7158 = 7158;
  localparam test_b1_S7159 = 7159;
  localparam test_b1_S7160 = 7160;
  localparam test_b1_S7161 = 7161;
  localparam test_b1_S7162 = 7162;
  localparam test_b1_S7163 = 7163;
  localparam test_b1_S7164 = 7164;
  localparam test_b1_S7165 = 7165;
  localparam test_b1_S7166 = 7166;
  localparam test_b1_S7167 = 7167;
  localparam test_b1_S7168 = 7168;
  localparam test_b1_S7169 = 7169;
  localparam test_b1_S7170 = 7170;
  localparam test_b1_S7171 = 7171;
  localparam test_b1_S7172 = 7172;
  localparam test_b1_S7173 = 7173;
  localparam test_b1_S7174 = 7174;
  localparam test_b1_S7175 = 7175;
  localparam test_b1_S7176 = 7176;
  localparam test_b1_S7177 = 7177;
  localparam test_b1_S7178 = 7178;
  localparam test_b1_S7179 = 7179;
  localparam test_b1_S7180 = 7180;
  localparam test_b1_S7181 = 7181;
  localparam test_b1_S7182 = 7182;
  localparam test_b1_S7183 = 7183;
  localparam test_b1_S7184 = 7184;
  localparam test_b1_S7185 = 7185;
  localparam test_b1_S7186 = 7186;
  localparam test_b1_S7187 = 7187;
  localparam test_b1_S7188 = 7188;
  localparam test_b1_S7189 = 7189;
  localparam test_b1_S7190 = 7190;
  localparam test_b1_S7191 = 7191;
  localparam test_b1_S7192 = 7192;
  localparam test_b1_S7193 = 7193;
  localparam test_b1_S7194 = 7194;
  localparam test_b1_S7195 = 7195;
  localparam test_b1_S7196 = 7196;
  localparam test_b1_S7197 = 7197;
  localparam test_b1_S7198 = 7198;
  localparam test_b1_S7199 = 7199;
  localparam test_b1_S7200 = 7200;
  localparam test_b1_S7201 = 7201;
  localparam test_b1_S7202 = 7202;
  localparam test_b1_S7203 = 7203;
  localparam test_b1_S7204 = 7204;
  localparam test_b1_S7205 = 7205;
  localparam test_b1_S7206 = 7206;
  localparam test_b1_S7207 = 7207;
  localparam test_b1_S7208 = 7208;
  localparam test_b1_S7209 = 7209;
  localparam test_b1_S7210 = 7210;
  localparam test_b1_S7211 = 7211;
  localparam test_b1_S7212 = 7212;
  localparam test_b1_S7213 = 7213;
  localparam test_b1_S7214 = 7214;
  localparam test_b1_S7215 = 7215;
  localparam test_b1_S7216 = 7216;
  localparam test_b1_S7217 = 7217;
  localparam test_b1_S7218 = 7218;
  localparam test_b1_S7219 = 7219;
  localparam test_b1_S7220 = 7220;
  localparam test_b1_S7221 = 7221;
  localparam test_b1_S7222 = 7222;
  localparam test_b1_S7223 = 7223;
  localparam test_b1_S7224 = 7224;
  localparam test_b1_S7225 = 7225;
  localparam test_b1_S7226 = 7226;
  localparam test_b1_S7227 = 7227;
  localparam test_b1_S7228 = 7228;
  localparam test_b1_S7229 = 7229;
  localparam test_b1_S7230 = 7230;
  localparam test_b1_S7231 = 7231;
  localparam test_b1_S7232 = 7232;
  localparam test_b1_S7233 = 7233;
  localparam test_b1_S7234 = 7234;
  localparam test_b1_S7235 = 7235;
  localparam test_b1_S7236 = 7236;
  localparam test_b1_S7237 = 7237;
  localparam test_b1_S7238 = 7238;
  localparam test_b1_S7239 = 7239;
  localparam test_b1_S7240 = 7240;
  localparam test_b1_S7241 = 7241;
  localparam test_b1_S7242 = 7242;
  localparam test_b1_S7243 = 7243;
  localparam test_b1_S7244 = 7244;
  localparam test_b1_S7245 = 7245;
  localparam test_b1_S7246 = 7246;
  localparam test_b1_S7247 = 7247;
  localparam test_b1_S7248 = 7248;
  localparam test_b1_S7249 = 7249;
  localparam test_b1_S7250 = 7250;
  localparam test_b1_S7251 = 7251;
  localparam test_b1_S7252 = 7252;
  localparam test_b1_S7253 = 7253;
  localparam test_b1_S7254 = 7254;
  localparam test_b1_S7255 = 7255;
  localparam test_b1_S7256 = 7256;
  localparam test_b1_S7257 = 7257;
  localparam test_b1_S7258 = 7258;
  localparam test_b1_S7259 = 7259;
  localparam test_b1_S7260 = 7260;
  localparam test_b1_S7261 = 7261;
  localparam test_b1_S7262 = 7262;
  localparam test_b1_S7263 = 7263;
  localparam test_b1_S7264 = 7264;
  localparam test_b1_S7265 = 7265;
  localparam test_b1_S7266 = 7266;
  localparam test_b1_S7267 = 7267;
  localparam test_b1_S7268 = 7268;
  localparam test_b1_S7269 = 7269;
  localparam test_b1_S7270 = 7270;
  localparam test_b1_S7271 = 7271;
  localparam test_b1_S7272 = 7272;
  localparam test_b1_S7273 = 7273;
  localparam test_b1_S7274 = 7274;
  localparam test_b1_S7275 = 7275;
  localparam test_b1_S7276 = 7276;
  localparam test_b1_S7277 = 7277;
  localparam test_b1_S7278 = 7278;
  localparam test_b1_S7279 = 7279;
  localparam test_b1_S7280 = 7280;
  localparam test_b1_S7281 = 7281;
  localparam test_b1_S7282 = 7282;
  localparam test_b1_S7283 = 7283;
  localparam test_b1_S7284 = 7284;
  localparam test_b1_S7285 = 7285;
  localparam test_b1_S7286 = 7286;
  localparam test_b1_S7287 = 7287;
  localparam test_b1_S7288 = 7288;
  localparam test_b1_S7289 = 7289;
  localparam test_b1_S7290 = 7290;
  localparam test_b1_S7291 = 7291;
  localparam test_b1_S7292 = 7292;
  localparam test_b1_S7293 = 7293;
  localparam test_b1_S7294 = 7294;
  localparam test_b1_S7295 = 7295;
  localparam test_b1_S7296 = 7296;
  localparam test_b1_S7297 = 7297;
  localparam test_b1_S7298 = 7298;
  localparam test_b1_S7299 = 7299;
  localparam test_b1_S7300 = 7300;
  localparam test_b1_S7301 = 7301;
  localparam test_b1_S7302 = 7302;
  localparam test_b1_S7303 = 7303;
  localparam test_b1_S7304 = 7304;
  localparam test_b1_S7305 = 7305;
  localparam test_b1_S7306 = 7306;
  localparam test_b1_S7307 = 7307;
  localparam test_b1_S7308 = 7308;
  localparam test_b1_S7309 = 7309;
  localparam test_b1_S7310 = 7310;
  localparam test_b1_S7311 = 7311;
  localparam test_b1_S7312 = 7312;
  localparam test_b1_S7313 = 7313;
  localparam test_b1_S7314 = 7314;
  localparam test_b1_S7315 = 7315;
  localparam test_b1_S7316 = 7316;
  localparam test_b1_S7317 = 7317;
  localparam test_b1_S7318 = 7318;
  localparam test_b1_S7319 = 7319;
  localparam test_b1_S7320 = 7320;
  localparam test_b1_S7321 = 7321;
  localparam test_b1_S7322 = 7322;
  localparam test_b1_S7323 = 7323;
  localparam test_b1_S7324 = 7324;
  localparam test_b1_S7325 = 7325;
  localparam test_b1_S7326 = 7326;
  localparam test_b1_S7327 = 7327;
  localparam test_b1_S7328 = 7328;
  localparam test_b1_S7329 = 7329;
  localparam test_b1_S7330 = 7330;
  localparam test_b1_S7331 = 7331;
  localparam test_b1_S7332 = 7332;
  localparam test_b1_S7333 = 7333;
  localparam test_b1_S7334 = 7334;
  localparam test_b1_S7335 = 7335;
  localparam test_b1_S7336 = 7336;
  localparam test_b1_S7337 = 7337;
  localparam test_b1_S7338 = 7338;
  localparam test_b1_S7339 = 7339;
  localparam test_b1_S7340 = 7340;
  localparam test_b1_S7341 = 7341;
  localparam test_b1_S7342 = 7342;
  localparam test_b1_S7343 = 7343;
  localparam test_b1_S7344 = 7344;
  localparam test_b1_S7345 = 7345;
  localparam test_b1_S7346 = 7346;
  localparam test_b1_S7347 = 7347;
  localparam test_b1_S7348 = 7348;
  localparam test_b1_S7349 = 7349;
  localparam test_b1_S7350 = 7350;
  localparam test_b1_S7351 = 7351;
  localparam test_b1_S7352 = 7352;
  localparam test_b1_S7353 = 7353;
  localparam test_b1_S7354 = 7354;
  localparam test_b1_S7355 = 7355;
  localparam test_b1_S7356 = 7356;
  localparam test_b1_S7357 = 7357;
  localparam test_b1_S7358 = 7358;
  localparam test_b1_S7359 = 7359;
  localparam test_b1_S7360 = 7360;
  localparam test_b1_S7361 = 7361;
  localparam test_b1_S7362 = 7362;
  localparam test_b1_S7363 = 7363;
  localparam test_b1_S7364 = 7364;
  localparam test_b1_S7365 = 7365;
  localparam test_b1_S7366 = 7366;
  localparam test_b1_S7367 = 7367;
  localparam test_b1_S7368 = 7368;
  localparam test_b1_S7369 = 7369;
  localparam test_b1_S7370 = 7370;
  localparam test_b1_S7371 = 7371;
  localparam test_b1_S7372 = 7372;
  localparam test_b1_S7373 = 7373;
  localparam test_b1_S7374 = 7374;
  localparam test_b1_S7375 = 7375;
  localparam test_b1_S7376 = 7376;
  localparam test_b1_S7377 = 7377;
  localparam test_b1_S7378 = 7378;
  localparam test_b1_S7379 = 7379;
  localparam test_b1_S7380 = 7380;
  localparam test_b1_S7381 = 7381;
  localparam test_b1_S7382 = 7382;
  localparam test_b1_S7383 = 7383;
  localparam test_b1_S7384 = 7384;
  localparam test_b1_S7385 = 7385;
  localparam test_b1_S7386 = 7386;
  localparam test_b1_S7387 = 7387;
  localparam test_b1_S7388 = 7388;
  localparam test_b1_S7389 = 7389;
  localparam test_b1_S7390 = 7390;
  localparam test_b1_S7391 = 7391;
  localparam test_b1_S7392 = 7392;
  localparam test_b1_S7393 = 7393;
  localparam test_b1_S7394 = 7394;
  localparam test_b1_S7395 = 7395;
  localparam test_b1_S7396 = 7396;
  localparam test_b1_S7397 = 7397;
  localparam test_b1_S7398 = 7398;
  localparam test_b1_S7399 = 7399;
  localparam test_b1_S7400 = 7400;
  localparam test_b1_S7401 = 7401;
  localparam test_b1_S7402 = 7402;
  localparam test_b1_S7403 = 7403;
  localparam test_b1_S7404 = 7404;
  localparam test_b1_S7405 = 7405;
  localparam test_b1_S7406 = 7406;
  localparam test_b1_S7407 = 7407;
  localparam test_b1_S7408 = 7408;
  localparam test_b1_S7409 = 7409;
  localparam test_b1_S7410 = 7410;
  localparam test_b1_S7411 = 7411;
  localparam test_b1_S7412 = 7412;
  localparam test_b1_S7413 = 7413;
  localparam test_b1_S7414 = 7414;
  localparam test_b1_S7415 = 7415;
  localparam test_b1_S7416 = 7416;
  localparam test_b1_S7417 = 7417;
  localparam test_b1_S7418 = 7418;
  localparam test_b1_S7419 = 7419;
  localparam test_b1_S7420 = 7420;
  localparam test_b1_S7421 = 7421;
  localparam test_b1_S7422 = 7422;
  localparam test_b1_S7423 = 7423;
  localparam test_b1_S7424 = 7424;
  localparam test_b1_S7425 = 7425;
  localparam test_b1_S7426 = 7426;
  localparam test_b1_S7427 = 7427;
  localparam test_b1_S7428 = 7428;
  localparam test_b1_S7429 = 7429;
  localparam test_b1_S7430 = 7430;
  localparam test_b1_S7431 = 7431;
  localparam test_b1_S7432 = 7432;
  localparam test_b1_S7433 = 7433;
  localparam test_b1_S7434 = 7434;
  localparam test_b1_S7435 = 7435;
  localparam test_b1_S7436 = 7436;
  localparam test_b1_S7437 = 7437;
  localparam test_b1_S7438 = 7438;
  localparam test_b1_S7439 = 7439;
  localparam test_b1_S7440 = 7440;
  localparam test_b1_S7441 = 7441;
  localparam test_b1_S7442 = 7442;
  localparam test_b1_S7443 = 7443;
  localparam test_b1_S7444 = 7444;
  localparam test_b1_S7445 = 7445;
  localparam test_b1_S7446 = 7446;
  localparam test_b1_S7447 = 7447;
  localparam test_b1_S7448 = 7448;
  localparam test_b1_S7449 = 7449;
  localparam test_b1_S7450 = 7450;
  localparam test_b1_S7451 = 7451;
  localparam test_b1_S7452 = 7452;
  localparam test_b1_S7453 = 7453;
  localparam test_b1_S7454 = 7454;
  localparam test_b1_S7455 = 7455;
  localparam test_b1_S7456 = 7456;
  localparam test_b1_S7457 = 7457;
  localparam test_b1_S7458 = 7458;
  localparam test_b1_S7459 = 7459;
  localparam test_b1_S7460 = 7460;
  localparam test_b1_S7461 = 7461;
  localparam test_b1_S7462 = 7462;
  localparam test_b1_S7463 = 7463;
  localparam test_b1_S7464 = 7464;
  localparam test_b1_S7465 = 7465;
  localparam test_b1_S7466 = 7466;
  localparam test_b1_S7467 = 7467;
  localparam test_b1_S7468 = 7468;
  localparam test_b1_S7469 = 7469;
  localparam test_b1_S7470 = 7470;
  localparam test_b1_S7471 = 7471;
  localparam test_b1_S7472 = 7472;
  localparam test_b1_S7473 = 7473;
  localparam test_b1_S7474 = 7474;
  localparam test_b1_S7475 = 7475;
  localparam test_b1_S7476 = 7476;
  localparam test_b1_S7477 = 7477;
  localparam test_b1_S7478 = 7478;
  localparam test_b1_S7479 = 7479;
  localparam test_b1_S7480 = 7480;
  localparam test_b1_S7481 = 7481;
  localparam test_b1_S7482 = 7482;
  localparam test_b1_S7483 = 7483;
  localparam test_b1_S7484 = 7484;
  localparam test_b1_S7485 = 7485;
  localparam test_b1_S7486 = 7486;
  localparam test_b1_S7487 = 7487;
  localparam test_b1_S7488 = 7488;
  localparam test_b1_S7489 = 7489;
  localparam test_b1_S7490 = 7490;
  localparam test_b1_S7491 = 7491;
  localparam test_b1_S7492 = 7492;
  localparam test_b1_S7493 = 7493;
  localparam test_b1_S7494 = 7494;
  localparam test_b1_S7495 = 7495;
  localparam test_b1_S7496 = 7496;
  localparam test_b1_S7497 = 7497;
  localparam test_b1_S7498 = 7498;
  localparam test_b1_S7499 = 7499;
  localparam test_b1_S7500 = 7500;
  localparam test_b1_S7501 = 7501;
  localparam test_b1_S7502 = 7502;
  localparam test_b1_S7503 = 7503;
  localparam test_b1_S7504 = 7504;
  localparam test_b1_S7505 = 7505;
  localparam test_b1_S7506 = 7506;
  localparam test_b1_S7507 = 7507;
  localparam test_b1_S7508 = 7508;
  localparam test_b1_S7509 = 7509;
  localparam test_b1_S7510 = 7510;
  localparam test_b1_S7511 = 7511;
  localparam test_b1_S7512 = 7512;
  localparam test_b1_S7513 = 7513;
  localparam test_b1_S7514 = 7514;
  localparam test_b1_S7515 = 7515;
  localparam test_b1_S7516 = 7516;
  localparam test_b1_S7517 = 7517;
  localparam test_b1_S7518 = 7518;
  localparam test_b1_S7519 = 7519;
  localparam test_b1_S7520 = 7520;
  localparam test_b1_S7521 = 7521;
  localparam test_b1_S7522 = 7522;
  localparam test_b1_S7523 = 7523;
  localparam test_b1_S7524 = 7524;
  localparam test_b1_S7525 = 7525;
  localparam test_b1_S7526 = 7526;
  localparam test_b1_S7527 = 7527;
  localparam test_b1_S7528 = 7528;
  localparam test_b1_S7529 = 7529;
  localparam test_b1_S7530 = 7530;
  localparam test_b1_S7531 = 7531;
  localparam test_b1_S7532 = 7532;
  localparam test_b1_S7533 = 7533;
  localparam test_b1_S7534 = 7534;
  localparam test_b1_S7535 = 7535;
  localparam test_b1_S7536 = 7536;
  localparam test_b1_S7537 = 7537;
  localparam test_b1_S7538 = 7538;
  localparam test_b1_S7539 = 7539;
  localparam test_b1_S7540 = 7540;
  localparam test_b1_S7541 = 7541;
  localparam test_b1_S7542 = 7542;
  localparam test_b1_S7543 = 7543;
  localparam test_b1_S7544 = 7544;
  localparam test_b1_S7545 = 7545;
  localparam test_b1_S7546 = 7546;
  localparam test_b1_S7547 = 7547;
  localparam test_b1_S7548 = 7548;
  localparam test_b1_S7549 = 7549;
  localparam test_b1_S7550 = 7550;
  localparam test_b1_S7551 = 7551;
  localparam test_b1_S7552 = 7552;
  localparam test_b1_S7553 = 7553;
  localparam test_b1_S7554 = 7554;
  localparam test_b1_S7555 = 7555;
  localparam test_b1_S7556 = 7556;
  localparam test_b1_S7557 = 7557;
  localparam test_b1_S7558 = 7558;
  localparam test_b1_S7559 = 7559;
  localparam test_b1_S7560 = 7560;
  localparam test_b1_S7561 = 7561;
  localparam test_b1_S7562 = 7562;
  localparam test_b1_S7563 = 7563;
  localparam test_b1_S7564 = 7564;
  localparam test_b1_S7565 = 7565;
  localparam test_b1_S7566 = 7566;
  localparam test_b1_S7567 = 7567;
  localparam test_b1_S7568 = 7568;
  localparam test_b1_S7569 = 7569;
  localparam test_b1_S7570 = 7570;
  localparam test_b1_S7571 = 7571;
  localparam test_b1_S7572 = 7572;
  localparam test_b1_S7573 = 7573;
  localparam test_b1_S7574 = 7574;
  localparam test_b1_S7575 = 7575;
  localparam test_b1_S7576 = 7576;
  localparam test_b1_S7577 = 7577;
  localparam test_b1_S7578 = 7578;
  localparam test_b1_S7579 = 7579;
  localparam test_b1_S7580 = 7580;
  localparam test_b1_S7581 = 7581;
  localparam test_b1_S7582 = 7582;
  localparam test_b1_S7583 = 7583;
  localparam test_b1_S7584 = 7584;
  localparam test_b1_S7585 = 7585;
  localparam test_b1_S7586 = 7586;
  localparam test_b1_S7587 = 7587;
  localparam test_b1_S7588 = 7588;
  localparam test_b1_S7589 = 7589;
  localparam test_b1_S7590 = 7590;
  localparam test_b1_S7591 = 7591;
  localparam test_b1_S7592 = 7592;
  localparam test_b1_S7593 = 7593;
  localparam test_b1_S7594 = 7594;
  localparam test_b1_S7595 = 7595;
  localparam test_b1_S7596 = 7596;
  localparam test_b1_S7597 = 7597;
  localparam test_b1_S7598 = 7598;
  localparam test_b1_S7599 = 7599;
  localparam test_b1_S7600 = 7600;
  localparam test_b1_S7601 = 7601;
  localparam test_b1_S7602 = 7602;
  localparam test_b1_S7603 = 7603;
  localparam test_b1_S7604 = 7604;
  localparam test_b1_S7605 = 7605;
  localparam test_b1_S7606 = 7606;
  localparam test_b1_S7607 = 7607;
  localparam test_b1_S7608 = 7608;
  localparam test_b1_S7609 = 7609;
  localparam test_b1_S7610 = 7610;
  localparam test_b1_S7611 = 7611;
  localparam test_b1_S7612 = 7612;
  localparam test_b1_S7613 = 7613;
  localparam test_b1_S7614 = 7614;
  localparam test_b1_S7615 = 7615;
  localparam test_b1_S7616 = 7616;
  localparam test_b1_S7617 = 7617;
  localparam test_b1_S7618 = 7618;
  localparam test_b1_S7619 = 7619;
  localparam test_b1_S7620 = 7620;
  localparam test_b1_S7621 = 7621;
  localparam test_b1_S7622 = 7622;
  localparam test_b1_S7623 = 7623;
  localparam test_b1_S7624 = 7624;
  localparam test_b1_S7625 = 7625;
  localparam test_b1_S7626 = 7626;
  localparam test_b1_S7627 = 7627;
  localparam test_b1_S7628 = 7628;
  localparam test_b1_S7629 = 7629;
  localparam test_b1_S7630 = 7630;
  localparam test_b1_S7631 = 7631;
  localparam test_b1_S7632 = 7632;
  localparam test_b1_S7633 = 7633;
  localparam test_b1_S7634 = 7634;
  localparam test_b1_S7635 = 7635;
  localparam test_b1_S7636 = 7636;
  localparam test_b1_S7637 = 7637;
  localparam test_b1_S7638 = 7638;
  localparam test_b1_S7639 = 7639;
  localparam test_b1_S7640 = 7640;
  localparam test_b1_S7641 = 7641;
  localparam test_b1_S7642 = 7642;
  localparam test_b1_S7643 = 7643;
  localparam test_b1_S7644 = 7644;
  localparam test_b1_S7645 = 7645;
  localparam test_b1_S7646 = 7646;
  localparam test_b1_S7647 = 7647;
  localparam test_b1_S7648 = 7648;
  localparam test_b1_S7649 = 7649;
  localparam test_b1_S7650 = 7650;
  localparam test_b1_S7651 = 7651;
  localparam test_b1_S7652 = 7652;
  localparam test_b1_S7653 = 7653;
  localparam test_b1_S7654 = 7654;
  localparam test_b1_S7655 = 7655;
  localparam test_b1_S7656 = 7656;
  localparam test_b1_S7657 = 7657;
  localparam test_b1_S7658 = 7658;
  localparam test_b1_S7659 = 7659;
  localparam test_b1_S7660 = 7660;
  localparam test_b1_S7661 = 7661;
  localparam test_b1_S7662 = 7662;
  localparam test_b1_S7663 = 7663;
  localparam test_b1_S7664 = 7664;
  localparam test_b1_S7665 = 7665;
  localparam test_b1_S7666 = 7666;
  localparam test_b1_S7667 = 7667;
  localparam test_b1_S7668 = 7668;
  localparam test_b1_S7669 = 7669;
  localparam test_b1_S7670 = 7670;
  localparam test_b1_S7671 = 7671;
  localparam test_b1_S7672 = 7672;
  localparam test_b1_S7673 = 7673;
  localparam test_b1_S7674 = 7674;
  localparam test_b1_S7675 = 7675;
  localparam test_b1_S7676 = 7676;
  localparam test_b1_S7677 = 7677;
  localparam test_b1_S7678 = 7678;
  localparam test_b1_S7679 = 7679;
  localparam test_b1_S7680 = 7680;
  localparam test_b1_S7681 = 7681;
  localparam test_b1_S7682 = 7682;
  localparam test_b1_S7683 = 7683;
  localparam test_b1_S7684 = 7684;
  localparam test_b1_S7685 = 7685;
  localparam test_b1_S7686 = 7686;
  localparam test_b1_S7687 = 7687;
  localparam test_b1_S7688 = 7688;
  localparam test_b1_S7689 = 7689;
  localparam test_b1_S7690 = 7690;
  localparam test_b1_S7691 = 7691;
  localparam test_b1_S7692 = 7692;
  localparam test_b1_S7693 = 7693;
  localparam test_b1_S7694 = 7694;
  localparam test_b1_S7695 = 7695;
  localparam test_b1_S7696 = 7696;
  localparam test_b1_S7697 = 7697;
  localparam test_b1_S7698 = 7698;
  localparam test_b1_S7699 = 7699;
  localparam test_b1_S7700 = 7700;
  localparam test_b1_S7701 = 7701;
  localparam test_b1_S7702 = 7702;
  localparam test_b1_S7703 = 7703;
  localparam test_b1_S7704 = 7704;
  localparam test_b1_S7705 = 7705;
  localparam test_b1_S7706 = 7706;
  localparam test_b1_S7707 = 7707;
  localparam test_b1_S7708 = 7708;
  localparam test_b1_S7709 = 7709;
  localparam test_b1_S7710 = 7710;
  localparam test_b1_S7711 = 7711;
  localparam test_b1_S7712 = 7712;
  localparam test_b1_S7713 = 7713;
  localparam test_b1_S7714 = 7714;
  localparam test_b1_S7715 = 7715;
  localparam test_b1_S7716 = 7716;
  localparam test_b1_S7717 = 7717;
  localparam test_b1_S7718 = 7718;
  localparam test_b1_S7719 = 7719;
  localparam test_b1_S7720 = 7720;
  localparam test_b1_S7721 = 7721;
  localparam test_b1_S7722 = 7722;
  localparam test_b1_S7723 = 7723;
  localparam test_b1_S7724 = 7724;
  localparam test_b1_S7725 = 7725;
  localparam test_b1_S7726 = 7726;
  localparam test_b1_S7727 = 7727;
  localparam test_b1_S7728 = 7728;
  localparam test_b1_S7729 = 7729;
  localparam test_b1_S7730 = 7730;
  localparam test_b1_S7731 = 7731;
  localparam test_b1_S7732 = 7732;
  localparam test_b1_S7733 = 7733;
  localparam test_b1_S7734 = 7734;
  localparam test_b1_S7735 = 7735;
  localparam test_b1_S7736 = 7736;
  localparam test_b1_S7737 = 7737;
  localparam test_b1_S7738 = 7738;
  localparam test_b1_S7739 = 7739;
  localparam test_b1_S7740 = 7740;
  localparam test_b1_S7741 = 7741;
  localparam test_b1_S7742 = 7742;
  localparam test_b1_S7743 = 7743;
  localparam test_b1_S7744 = 7744;
  localparam test_b1_S7745 = 7745;
  localparam test_b1_S7746 = 7746;
  localparam test_b1_S7747 = 7747;
  localparam test_b1_S7748 = 7748;
  localparam test_b1_S7749 = 7749;
  localparam test_b1_S7750 = 7750;
  localparam test_b1_S7751 = 7751;
  localparam test_b1_S7752 = 7752;
  localparam test_b1_S7753 = 7753;
  localparam test_b1_S7754 = 7754;
  localparam test_b1_S7755 = 7755;
  localparam test_b1_S7756 = 7756;
  localparam test_b1_S7757 = 7757;
  localparam test_b1_S7758 = 7758;
  localparam test_b1_S7759 = 7759;
  localparam test_b1_S7760 = 7760;
  localparam test_b1_S7761 = 7761;
  localparam test_b1_S7762 = 7762;
  localparam test_b1_S7763 = 7763;
  localparam test_b1_S7764 = 7764;
  localparam test_b1_S7765 = 7765;
  localparam test_b1_S7766 = 7766;
  localparam test_b1_S7767 = 7767;
  localparam test_b1_S7768 = 7768;
  localparam test_b1_S7769 = 7769;
  localparam test_b1_S7770 = 7770;
  localparam test_b1_S7771 = 7771;
  localparam test_b1_S7772 = 7772;
  localparam test_b1_S7773 = 7773;
  localparam test_b1_S7774 = 7774;
  localparam test_b1_S7775 = 7775;
  localparam test_b1_S7776 = 7776;
  localparam test_b1_S7777 = 7777;
  localparam test_b1_S7778 = 7778;
  localparam test_b1_S7779 = 7779;
  localparam test_b1_S7780 = 7780;
  localparam test_b1_S7781 = 7781;
  localparam test_b1_S7782 = 7782;
  localparam test_b1_S7783 = 7783;
  localparam test_b1_S7784 = 7784;
  localparam test_b1_S7785 = 7785;
  localparam test_b1_S7786 = 7786;
  localparam test_b1_S7787 = 7787;
  localparam test_b1_S7788 = 7788;
  localparam test_b1_S7789 = 7789;
  localparam test_b1_S7790 = 7790;
  localparam test_b1_S7791 = 7791;
  localparam test_b1_S7792 = 7792;
  localparam test_b1_S7793 = 7793;
  localparam test_b1_S7794 = 7794;
  localparam test_b1_S7795 = 7795;
  localparam test_b1_S7796 = 7796;
  localparam test_b1_S7797 = 7797;
  localparam test_b1_S7798 = 7798;
  localparam test_b1_S7799 = 7799;
  localparam test_b1_S7800 = 7800;
  localparam test_b1_S7801 = 7801;
  localparam test_b1_S7802 = 7802;
  localparam test_b1_S7803 = 7803;
  localparam test_b1_S7804 = 7804;
  localparam test_b1_S7805 = 7805;
  localparam test_b1_S7806 = 7806;
  localparam test_b1_S7807 = 7807;
  localparam test_b1_S7808 = 7808;
  localparam test_b1_S7809 = 7809;
  localparam test_b1_S7810 = 7810;
  localparam test_b1_S7811 = 7811;
  localparam test_b1_S7812 = 7812;
  localparam test_b1_S7813 = 7813;
  localparam test_b1_S7814 = 7814;
  localparam test_b1_S7815 = 7815;
  localparam test_b1_S7816 = 7816;
  localparam test_b1_S7817 = 7817;
  localparam test_b1_S7818 = 7818;
  localparam test_b1_S7819 = 7819;
  localparam test_b1_S7820 = 7820;
  localparam test_b1_S7821 = 7821;
  localparam test_b1_S7822 = 7822;
  localparam test_b1_S7823 = 7823;
  localparam test_b1_S7824 = 7824;
  localparam test_b1_S7825 = 7825;
  localparam test_b1_S7826 = 7826;
  localparam test_b1_S7827 = 7827;
  localparam test_b1_S7828 = 7828;
  localparam test_b1_S7829 = 7829;
  localparam test_b1_S7830 = 7830;
  localparam test_b1_S7831 = 7831;
  localparam test_b1_S7832 = 7832;
  localparam test_b1_S7833 = 7833;
  localparam test_b1_S7834 = 7834;
  localparam test_b1_S7835 = 7835;
  localparam test_b1_S7836 = 7836;
  localparam test_b1_S7837 = 7837;
  localparam test_b1_S7838 = 7838;
  localparam test_b1_S7839 = 7839;
  localparam test_b1_S7840 = 7840;
  localparam test_b1_S7841 = 7841;
  localparam test_b1_S7842 = 7842;
  localparam test_b1_S7843 = 7843;
  localparam test_b1_S7844 = 7844;
  localparam test_b1_S7845 = 7845;
  localparam test_b1_S7846 = 7846;
  localparam test_b1_S7847 = 7847;
  localparam test_b1_S7848 = 7848;
  localparam test_b1_S7849 = 7849;
  localparam test_b1_S7850 = 7850;
  localparam test_b1_S7851 = 7851;
  localparam test_b1_S7852 = 7852;
  localparam test_b1_S7853 = 7853;
  localparam test_b1_S7854 = 7854;
  localparam test_b1_S7855 = 7855;
  localparam test_b1_S7856 = 7856;
  localparam test_b1_S7857 = 7857;
  localparam test_b1_S7858 = 7858;
  localparam test_b1_S7859 = 7859;
  localparam test_b1_S7860 = 7860;
  localparam test_b1_S7861 = 7861;
  localparam test_b1_S7862 = 7862;
  localparam test_b1_S7863 = 7863;
  localparam test_b1_S7864 = 7864;
  localparam test_b1_S7865 = 7865;
  localparam test_b1_S7866 = 7866;
  localparam test_b1_S7867 = 7867;
  localparam test_b1_S7868 = 7868;
  localparam test_b1_S7869 = 7869;
  localparam test_b1_S7870 = 7870;
  localparam test_b1_S7871 = 7871;
  localparam test_b1_S7872 = 7872;
  localparam test_b1_S7873 = 7873;
  localparam test_b1_S7874 = 7874;
  localparam test_b1_S7875 = 7875;
  localparam test_b1_S7876 = 7876;
  localparam test_b1_S7877 = 7877;
  localparam test_b1_S7878 = 7878;
  localparam test_b1_S7879 = 7879;
  localparam test_b1_S7880 = 7880;
  localparam test_b1_S7881 = 7881;
  localparam test_b1_S7882 = 7882;
  localparam test_b1_S7883 = 7883;
  localparam test_b1_S7884 = 7884;
  localparam test_b1_S7885 = 7885;
  localparam test_b1_S7886 = 7886;
  localparam test_b1_S7887 = 7887;
  localparam test_b1_S7888 = 7888;
  localparam test_b1_S7889 = 7889;
  localparam test_b1_S7890 = 7890;
  localparam test_b1_S7891 = 7891;
  localparam test_b1_S7892 = 7892;
  localparam test_b1_S7893 = 7893;
  localparam test_b1_S7894 = 7894;
  localparam test_b1_S7895 = 7895;
  localparam test_b1_S7896 = 7896;
  localparam test_b1_S7897 = 7897;
  localparam test_b1_S7898 = 7898;
  localparam test_b1_S7899 = 7899;
  localparam test_b1_S7900 = 7900;
  localparam test_b1_S7901 = 7901;
  localparam test_b1_S7902 = 7902;
  localparam test_b1_S7903 = 7903;
  localparam test_b1_S7904 = 7904;
  localparam test_b1_S7905 = 7905;
  localparam test_b1_S7906 = 7906;
  localparam test_b1_S7907 = 7907;
  localparam test_b1_S7908 = 7908;
  localparam test_b1_S7909 = 7909;
  localparam test_b1_S7910 = 7910;
  localparam test_b1_S7911 = 7911;
  localparam test_b1_S7912 = 7912;
  localparam test_b1_S7913 = 7913;
  localparam test_b1_S7914 = 7914;
  localparam test_b1_S7915 = 7915;
  localparam test_b1_S7916 = 7916;
  localparam test_b1_S7917 = 7917;
  localparam test_b1_S7918 = 7918;
  localparam test_b1_S7919 = 7919;
  localparam test_b1_S7920 = 7920;
  localparam test_b1_S7921 = 7921;
  localparam test_b1_S7922 = 7922;
  localparam test_b1_S7923 = 7923;
  localparam test_b1_S7924 = 7924;
  localparam test_b1_S7925 = 7925;
  localparam test_b1_S7926 = 7926;
  localparam test_b1_S7927 = 7927;
  localparam test_b1_S7928 = 7928;
  localparam test_b1_S7929 = 7929;
  localparam test_b1_S7930 = 7930;
  localparam test_b1_S7931 = 7931;
  localparam test_b1_S7932 = 7932;
  localparam test_b1_S7933 = 7933;
  localparam test_b1_S7934 = 7934;
  localparam test_b1_S7935 = 7935;
  localparam test_b1_S7936 = 7936;
  localparam test_b1_S7937 = 7937;
  localparam test_b1_S7938 = 7938;
  localparam test_b1_S7939 = 7939;
  localparam test_b1_S7940 = 7940;
  localparam test_b1_S7941 = 7941;
  localparam test_b1_S7942 = 7942;
  localparam test_b1_S7943 = 7943;
  localparam test_b1_S7944 = 7944;
  localparam test_b1_S7945 = 7945;
  localparam test_b1_S7946 = 7946;
  localparam test_b1_S7947 = 7947;
  localparam test_b1_S7948 = 7948;
  localparam test_b1_S7949 = 7949;
  localparam test_b1_S7950 = 7950;
  localparam test_b1_S7951 = 7951;
  localparam test_b1_S7952 = 7952;
  localparam test_b1_S7953 = 7953;
  localparam test_b1_S7954 = 7954;
  localparam test_b1_S7955 = 7955;
  localparam test_b1_S7956 = 7956;
  localparam test_b1_S7957 = 7957;
  localparam test_b1_S7958 = 7958;
  localparam test_b1_S7959 = 7959;
  localparam test_b1_S7960 = 7960;
  localparam test_b1_S7961 = 7961;
  localparam test_b1_S7962 = 7962;
  localparam test_b1_S7963 = 7963;
  localparam test_b1_S7964 = 7964;
  localparam test_b1_S7965 = 7965;
  localparam test_b1_S7966 = 7966;
  localparam test_b1_S7967 = 7967;
  localparam test_b1_S7968 = 7968;
  localparam test_b1_S7969 = 7969;
  localparam test_b1_S7970 = 7970;
  localparam test_b1_S7971 = 7971;
  localparam test_b1_S7972 = 7972;
  localparam test_b1_S7973 = 7973;
  localparam test_b1_S7974 = 7974;
  localparam test_b1_S7975 = 7975;
  localparam test_b1_S7976 = 7976;
  localparam test_b1_S7977 = 7977;
  localparam test_b1_S7978 = 7978;
  localparam test_b1_S7979 = 7979;
  localparam test_b1_S7980 = 7980;
  localparam test_b1_S7981 = 7981;
  localparam test_b1_S7982 = 7982;
  localparam test_b1_S7983 = 7983;
  localparam test_b1_S7984 = 7984;
  localparam test_b1_S7985 = 7985;
  localparam test_b1_S7986 = 7986;
  localparam test_b1_S7987 = 7987;
  localparam test_b1_S7988 = 7988;
  localparam test_b1_S7989 = 7989;
  localparam test_b1_S7990 = 7990;
  localparam test_b1_S7991 = 7991;
  localparam test_b1_S7992 = 7992;
  localparam test_b1_S7993 = 7993;
  localparam test_b1_S7994 = 7994;
  localparam test_b1_S7995 = 7995;
  localparam test_b1_S7996 = 7996;
  localparam test_b1_S7997 = 7997;
  localparam test_b1_S7998 = 7998;
  localparam test_b1_S7999 = 7999;
  localparam test_b1_S8000 = 8000;
  localparam test_b1_S8001 = 8001;
  localparam test_b1_S8002 = 8002;
  localparam test_b1_S8003 = 8003;
  localparam test_b1_S8004 = 8004;
  localparam test_b1_S8005 = 8005;
  localparam test_b1_S8006 = 8006;
  localparam test_b1_S8007 = 8007;
  localparam test_b1_S8008 = 8008;
  localparam test_b1_S8009 = 8009;
  localparam test_b1_S8010 = 8010;
  localparam test_b1_S8011 = 8011;
  localparam test_b1_S8012 = 8012;
  localparam test_b1_S8013 = 8013;
  localparam test_b1_S8014 = 8014;
  localparam test_b1_S8015 = 8015;
  localparam test_b1_S8016 = 8016;
  localparam test_b1_S8017 = 8017;
  localparam test_b1_S8018 = 8018;
  localparam test_b1_S8019 = 8019;
  localparam test_b1_S8020 = 8020;
  localparam test_b1_S8021 = 8021;
  localparam test_b1_S8022 = 8022;
  localparam test_b1_S8023 = 8023;
  localparam test_b1_S8024 = 8024;
  localparam test_b1_S8025 = 8025;
  localparam test_b1_S8026 = 8026;
  localparam test_b1_S8027 = 8027;
  localparam test_b1_S8028 = 8028;
  localparam test_b1_S8029 = 8029;
  localparam test_b1_S8030 = 8030;
  localparam test_b1_S8031 = 8031;
  localparam test_b1_S8032 = 8032;
  localparam test_b1_S8033 = 8033;
  localparam test_b1_S8034 = 8034;
  localparam test_b1_S8035 = 8035;
  localparam test_b1_S8036 = 8036;
  localparam test_b1_S8037 = 8037;
  localparam test_b1_S8038 = 8038;
  localparam test_b1_S8039 = 8039;
  localparam test_b1_S8040 = 8040;
  localparam test_b1_S8041 = 8041;
  localparam test_b1_S8042 = 8042;
  localparam test_b1_S8043 = 8043;
  localparam test_b1_S8044 = 8044;
  localparam test_b1_S8045 = 8045;
  localparam test_b1_S8046 = 8046;
  localparam test_b1_S8047 = 8047;
  localparam test_b1_S8048 = 8048;
  localparam test_b1_S8049 = 8049;
  localparam test_b1_S8050 = 8050;
  localparam test_b1_S8051 = 8051;
  localparam test_b1_S8052 = 8052;
  localparam test_b1_S8053 = 8053;
  localparam test_b1_S8054 = 8054;
  localparam test_b1_S8055 = 8055;
  localparam test_b1_S8056 = 8056;
  localparam test_b1_S8057 = 8057;
  localparam test_b1_S8058 = 8058;
  localparam test_b1_S8059 = 8059;
  localparam test_b1_S8060 = 8060;
  localparam test_b1_S8061 = 8061;
  localparam test_b1_S8062 = 8062;
  localparam test_b1_S8063 = 8063;
  localparam test_b1_S8064 = 8064;
  localparam test_b1_S8065 = 8065;
  localparam test_b1_S8066 = 8066;
  localparam test_b1_S8067 = 8067;
  localparam test_b1_S8068 = 8068;
  localparam test_b1_S8069 = 8069;
  localparam test_b1_S8070 = 8070;
  localparam test_b1_S8071 = 8071;
  localparam test_b1_S8072 = 8072;
  localparam test_b1_S8073 = 8073;
  localparam test_b1_S8074 = 8074;
  localparam test_b1_S8075 = 8075;
  localparam test_b1_S8076 = 8076;
  localparam test_b1_S8077 = 8077;
  localparam test_b1_S8078 = 8078;
  localparam test_b1_S8079 = 8079;
  localparam test_b1_S8080 = 8080;
  localparam test_b1_S8081 = 8081;
  localparam test_b1_S8082 = 8082;
  localparam test_b1_S8083 = 8083;
  localparam test_b1_S8084 = 8084;
  localparam test_b1_S8085 = 8085;
  localparam test_b1_S8086 = 8086;
  localparam test_b1_S8087 = 8087;
  localparam test_b1_S8088 = 8088;
  localparam test_b1_S8089 = 8089;
  localparam test_b1_S8090 = 8090;
  localparam test_b1_S8091 = 8091;
  localparam test_b1_S8092 = 8092;
  localparam test_b1_S8093 = 8093;
  localparam test_b1_S8094 = 8094;
  localparam test_b1_S8095 = 8095;
  localparam test_b1_S8096 = 8096;
  localparam test_b1_S8097 = 8097;
  localparam test_b1_S8098 = 8098;
  localparam test_b1_S8099 = 8099;
  localparam test_b1_S8100 = 8100;
  localparam test_b1_S8101 = 8101;
  localparam test_b1_S8102 = 8102;
  localparam test_b1_S8103 = 8103;
  localparam test_b1_S8104 = 8104;
  localparam test_b1_S8105 = 8105;
  localparam test_b1_S8106 = 8106;
  localparam test_b1_S8107 = 8107;
  localparam test_b1_S8108 = 8108;
  localparam test_b1_S8109 = 8109;
  localparam test_b1_S8110 = 8110;
  localparam test_b1_S8111 = 8111;
  localparam test_b1_S8112 = 8112;
  localparam test_b1_S8113 = 8113;
  localparam test_b1_S8114 = 8114;
  localparam test_b1_S8115 = 8115;
  localparam test_b1_S8116 = 8116;
  localparam test_b1_S8117 = 8117;
  localparam test_b1_S8118 = 8118;
  localparam test_b1_S8119 = 8119;
  localparam test_b1_S8120 = 8120;
  localparam test_b1_S8121 = 8121;
  localparam test_b1_S8122 = 8122;
  localparam test_b1_S8123 = 8123;
  localparam test_b1_S8124 = 8124;
  localparam test_b1_S8125 = 8125;
  localparam test_b1_S8126 = 8126;
  localparam test_b1_S8127 = 8127;
  localparam test_b1_S8128 = 8128;
  localparam test_b1_S8129 = 8129;
  localparam test_b1_S8130 = 8130;
  localparam test_b1_S8131 = 8131;
  localparam test_b1_S8132 = 8132;
  localparam test_b1_S8133 = 8133;
  localparam test_b1_S8134 = 8134;
  localparam test_b1_S8135 = 8135;
  localparam test_b1_S8136 = 8136;
  localparam test_b1_S8137 = 8137;
  localparam test_b1_S8138 = 8138;
  localparam test_b1_S8139 = 8139;
  localparam test_b1_S8140 = 8140;
  localparam test_b1_S8141 = 8141;
  localparam test_b1_S8142 = 8142;
  localparam test_b1_S8143 = 8143;
  localparam test_b1_S8144 = 8144;
  localparam test_b1_S8145 = 8145;
  localparam test_b1_S8146 = 8146;
  localparam test_b1_S8147 = 8147;
  localparam test_b1_S8148 = 8148;
  localparam test_b1_S8149 = 8149;
  localparam test_b1_S8150 = 8150;
  localparam test_b1_S8151 = 8151;
  localparam test_b1_S8152 = 8152;
  localparam test_b1_S8153 = 8153;
  localparam test_b1_S8154 = 8154;
  localparam test_b1_S8155 = 8155;
  localparam test_b1_S8156 = 8156;
  localparam test_b1_S8157 = 8157;
  localparam test_b1_S8158 = 8158;
  localparam test_b1_S8159 = 8159;
  localparam test_b1_S8160 = 8160;
  localparam test_b1_S8161 = 8161;
  localparam test_b1_S8162 = 8162;
  localparam test_b1_S8163 = 8163;
  localparam test_b1_S8164 = 8164;
  localparam test_b1_S8165 = 8165;
  localparam test_b1_S8166 = 8166;
  localparam test_b1_S8167 = 8167;
  localparam test_b1_S8168 = 8168;
  localparam test_b1_S8169 = 8169;
  localparam test_b1_S8170 = 8170;
  localparam test_b1_S8171 = 8171;
  localparam test_b1_S8172 = 8172;
  localparam test_b1_S8173 = 8173;
  localparam test_b1_S8174 = 8174;
  localparam test_b1_S8175 = 8175;
  localparam test_b1_S8176 = 8176;
  localparam test_b1_S8177 = 8177;
  localparam test_b1_S8178 = 8178;
  localparam test_b1_S8179 = 8179;
  localparam test_b1_S8180 = 8180;
  localparam test_b1_S8181 = 8181;
  localparam test_b1_S8182 = 8182;
  localparam test_b1_S8183 = 8183;
  localparam test_b1_S8184 = 8184;
  localparam test_b1_S8185 = 8185;
  localparam test_b1_S8186 = 8186;
  localparam test_b1_S8187 = 8187;
  localparam test_b1_S8188 = 8188;
  localparam test_b1_S8189 = 8189;
  localparam test_b1_S8190 = 8190;
  localparam test_b1_S8191 = 8191;
  localparam test_b1_S8192 = 8192;
  localparam test_b1_S8193 = 8193;
  localparam test_b1_S8194 = 8194;
  localparam test_b1_S8195 = 8195;
  localparam test_b1_S8196 = 8196;
  localparam test_b1_S8197 = 8197;
  localparam test_b1_S8198 = 8198;
  localparam test_b1_S8199 = 8199;
  localparam test_b1_S8200 = 8200;
  localparam test_b1_S8201 = 8201;
  localparam test_b1_S8202 = 8202;
  localparam test_b1_S8203 = 8203;
  localparam test_b1_S8204 = 8204;
  localparam test_b1_S8205 = 8205;
  localparam test_b1_S8206 = 8206;
  localparam test_b1_S8207 = 8207;
  localparam test_b1_S8208 = 8208;
  localparam test_b1_S8209 = 8209;
  localparam test_b1_S8210 = 8210;
  localparam test_b1_S8211 = 8211;
  localparam test_b1_S8212 = 8212;
  localparam test_b1_S8213 = 8213;
  localparam test_b1_S8214 = 8214;
  localparam test_b1_S8215 = 8215;
  localparam test_b1_S8216 = 8216;
  localparam test_b1_S8217 = 8217;
  localparam test_b1_S8218 = 8218;
  localparam test_b1_S8219 = 8219;
  localparam test_b1_S8220 = 8220;
  localparam test_b1_S8221 = 8221;
  localparam test_b1_S8222 = 8222;
  localparam test_b1_S8223 = 8223;
  localparam test_b1_S8224 = 8224;
  localparam test_b1_S8225 = 8225;
  localparam test_b1_S8226 = 8226;
  localparam test_b1_S8227 = 8227;
  localparam test_b1_S8228 = 8228;
  localparam test_b1_S8229 = 8229;
  localparam test_b1_S8230 = 8230;
  localparam test_b1_S8231 = 8231;
  localparam test_b1_S8232 = 8232;
  localparam test_b1_S8233 = 8233;
  localparam test_b1_S8234 = 8234;
  localparam test_b1_S8235 = 8235;
  localparam test_b1_S8236 = 8236;
  localparam test_b1_S8237 = 8237;
  localparam test_b1_S8238 = 8238;
  localparam test_b1_S8239 = 8239;
  localparam test_b1_S8240 = 8240;
  localparam test_b1_S8241 = 8241;
  localparam test_b1_S8242 = 8242;
  localparam test_b1_S8243 = 8243;
  localparam test_b1_S8244 = 8244;
  localparam test_b1_S8245 = 8245;
  localparam test_b1_S8246 = 8246;
  localparam test_b1_S8247 = 8247;
  localparam test_b1_S8248 = 8248;
  localparam test_b1_S8249 = 8249;
  localparam test_b1_S8250 = 8250;
  localparam test_b1_S8251 = 8251;
  localparam test_b1_S8252 = 8252;
  localparam test_b1_S8253 = 8253;
  localparam test_b1_S8254 = 8254;
  localparam test_b1_S8255 = 8255;
  localparam test_b1_S8256 = 8256;
  localparam test_b1_S8257 = 8257;
  localparam test_b1_S8258 = 8258;
  localparam test_b1_S8259 = 8259;
  localparam test_b1_S8260 = 8260;
  localparam test_b1_S8261 = 8261;
  localparam test_b1_S8262 = 8262;
  localparam test_b1_S8263 = 8263;
  localparam test_b1_S8264 = 8264;
  localparam test_b1_S8265 = 8265;
  localparam test_b1_S8266 = 8266;
  localparam test_b1_S8267 = 8267;
  localparam test_b1_S8268 = 8268;
  localparam test_b1_S8269 = 8269;
  localparam test_b1_S8270 = 8270;
  localparam test_b1_S8271 = 8271;
  localparam test_b1_S8272 = 8272;
  localparam test_b1_S8273 = 8273;
  localparam test_b1_S8274 = 8274;
  localparam test_b1_S8275 = 8275;
  localparam test_b1_S8276 = 8276;
  localparam test_b1_S8277 = 8277;
  localparam test_b1_S8278 = 8278;
  localparam test_b1_S8279 = 8279;
  localparam test_b1_S8280 = 8280;
  localparam test_b1_S8281 = 8281;
  localparam test_b1_S8282 = 8282;
  localparam test_b1_S8283 = 8283;
  localparam test_b1_S8284 = 8284;
  localparam test_b1_S8285 = 8285;
  localparam test_b1_S8286 = 8286;
  localparam test_b1_S8287 = 8287;
  localparam test_b1_S8288 = 8288;
  localparam test_b1_S8289 = 8289;
  localparam test_b1_S8290 = 8290;
  localparam test_b1_S8291 = 8291;
  localparam test_b1_S8292 = 8292;
  localparam test_b1_S8293 = 8293;
  localparam test_b1_S8294 = 8294;
  localparam test_b1_S8295 = 8295;
  localparam test_b1_S8296 = 8296;
  localparam test_b1_S8297 = 8297;
  localparam test_b1_S8298 = 8298;
  localparam test_b1_S8299 = 8299;
  localparam test_b1_S8300 = 8300;
  localparam test_b1_S8301 = 8301;
  localparam test_b1_S8302 = 8302;
  localparam test_b1_S8303 = 8303;
  localparam test_b1_S8304 = 8304;
  localparam test_b1_S8305 = 8305;
  localparam test_b1_S8306 = 8306;
  localparam test_b1_S8307 = 8307;
  localparam test_b1_S8308 = 8308;
  localparam test_b1_S8309 = 8309;
  localparam test_b1_S8310 = 8310;
  localparam test_b1_S8311 = 8311;
  localparam test_b1_S8312 = 8312;
  localparam test_b1_S8313 = 8313;
  localparam test_b1_S8314 = 8314;
  localparam test_b1_S8315 = 8315;
  localparam test_b1_S8316 = 8316;
  localparam test_b1_S8317 = 8317;
  localparam test_b1_S8318 = 8318;
  localparam test_b1_S8319 = 8319;
  localparam test_b1_S8320 = 8320;
  localparam test_b1_S8321 = 8321;
  localparam test_b1_S8322 = 8322;
  localparam test_b1_S8323 = 8323;
  localparam test_b1_S8324 = 8324;
  localparam test_b1_S8325 = 8325;
  localparam test_b1_S8326 = 8326;
  localparam test_b1_S8327 = 8327;
  localparam test_b1_S8328 = 8328;
  localparam test_b1_S8329 = 8329;
  localparam test_b1_S8330 = 8330;
  localparam test_b1_S8331 = 8331;
  localparam test_b1_S8332 = 8332;
  localparam test_b1_S8333 = 8333;
  localparam test_b1_S8334 = 8334;
  localparam test_b1_S8335 = 8335;
  localparam test_b1_S8336 = 8336;
  localparam test_b1_S8337 = 8337;
  localparam test_b1_S8338 = 8338;
  localparam test_b1_S8339 = 8339;
  localparam test_b1_S8340 = 8340;
  localparam test_b1_S8341 = 8341;
  localparam test_b1_S8342 = 8342;
  localparam test_b1_S8343 = 8343;
  localparam test_b1_S8344 = 8344;
  localparam test_b1_S8345 = 8345;
  localparam test_b1_S8346 = 8346;
  localparam test_b1_S8347 = 8347;
  localparam test_b1_S8348 = 8348;
  localparam test_b1_S8349 = 8349;
  localparam test_b1_S8350 = 8350;
  localparam test_b1_S8351 = 8351;
  localparam test_b1_S8352 = 8352;
  localparam test_b1_S8353 = 8353;
  localparam test_b1_S8354 = 8354;
  localparam test_b1_S8355 = 8355;
  localparam test_b1_S8356 = 8356;
  localparam test_b1_S8357 = 8357;
  localparam test_b1_S8358 = 8358;
  localparam test_b1_S8359 = 8359;
  localparam test_b1_S8360 = 8360;
  localparam test_b1_S8361 = 8361;
  localparam test_b1_S8362 = 8362;
  localparam test_b1_S8363 = 8363;
  localparam test_b1_S8364 = 8364;
  localparam test_b1_S8365 = 8365;
  localparam test_b1_S8366 = 8366;
  localparam test_b1_S8367 = 8367;
  localparam test_b1_S8368 = 8368;
  localparam test_b1_S8369 = 8369;
  localparam test_b1_S8370 = 8370;
  localparam test_b1_S8371 = 8371;
  localparam test_b1_S8372 = 8372;
  localparam test_b1_S8373 = 8373;
  localparam test_b1_S8374 = 8374;
  localparam test_b1_S8375 = 8375;
  localparam test_b1_S8376 = 8376;
  localparam test_b1_S8377 = 8377;
  localparam test_b1_S8378 = 8378;
  localparam test_b1_S8379 = 8379;
  localparam test_b1_S8380 = 8380;
  localparam test_b1_S8381 = 8381;
  localparam test_b1_S8382 = 8382;
  localparam test_b1_S8383 = 8383;
  localparam test_b1_S8384 = 8384;
  localparam test_b1_S8385 = 8385;
  localparam test_b1_S8386 = 8386;
  localparam test_b1_S8387 = 8387;
  localparam test_b1_S8388 = 8388;
  localparam test_b1_S8389 = 8389;
  localparam test_b1_S8390 = 8390;
  localparam test_b1_S8391 = 8391;
  localparam test_b1_S8392 = 8392;
  localparam test_b1_S8393 = 8393;
  localparam test_b1_S8394 = 8394;
  localparam test_b1_S8395 = 8395;
  localparam test_b1_S8396 = 8396;
  localparam test_b1_S8397 = 8397;
  localparam test_b1_S8398 = 8398;
  localparam test_b1_S8399 = 8399;
  localparam test_b1_S8400 = 8400;
  localparam test_b1_S8401 = 8401;
  localparam test_b1_S8402 = 8402;
  localparam test_b1_S8403 = 8403;
  localparam test_b1_S8404 = 8404;
  localparam test_b1_S8405 = 8405;
  localparam test_b1_S8406 = 8406;
  localparam test_b1_S8407 = 8407;
  localparam test_b1_S8408 = 8408;
  localparam test_b1_S8409 = 8409;
  localparam test_b1_S8410 = 8410;
  localparam test_b1_S8411 = 8411;
  localparam test_b1_S8412 = 8412;
  localparam test_b1_S8413 = 8413;
  localparam test_b1_S8414 = 8414;
  localparam test_b1_S8415 = 8415;
  localparam test_b1_S8416 = 8416;
  localparam test_b1_S8417 = 8417;
  localparam test_b1_S8418 = 8418;
  localparam test_b1_S8419 = 8419;
  localparam test_b1_S8420 = 8420;
  localparam test_b1_S8421 = 8421;
  localparam test_b1_S8422 = 8422;
  localparam test_b1_S8423 = 8423;
  localparam test_b1_S8424 = 8424;
  localparam test_b1_S8425 = 8425;
  localparam test_b1_S8426 = 8426;
  localparam test_b1_S8427 = 8427;
  localparam test_b1_S8428 = 8428;
  localparam test_b1_S8429 = 8429;
  localparam test_b1_S8430 = 8430;
  localparam test_b1_S8431 = 8431;
  localparam test_b1_S8432 = 8432;
  localparam test_b1_S8433 = 8433;
  localparam test_b1_S8434 = 8434;
  localparam test_b1_S8435 = 8435;
  localparam test_b1_S8436 = 8436;
  localparam test_b1_S8437 = 8437;
  localparam test_b1_S8438 = 8438;
  localparam test_b1_S8439 = 8439;
  localparam test_b1_S8440 = 8440;
  localparam test_b1_S8441 = 8441;
  localparam test_b1_S8442 = 8442;
  localparam test_b1_S8443 = 8443;
  localparam test_b1_S8444 = 8444;
  localparam test_b1_S8445 = 8445;
  localparam test_b1_S8446 = 8446;
  localparam test_b1_S8447 = 8447;
  localparam test_b1_S8448 = 8448;
  localparam test_b1_S8449 = 8449;
  localparam test_b1_S8450 = 8450;
  localparam test_b1_S8451 = 8451;
  localparam test_b1_S8452 = 8452;
  localparam test_b1_S8453 = 8453;
  localparam test_b1_S8454 = 8454;
  localparam test_b1_S8455 = 8455;
  localparam test_b1_S8456 = 8456;
  localparam test_b1_S8457 = 8457;
  localparam test_b1_S8458 = 8458;
  localparam test_b1_S8459 = 8459;
  localparam test_b1_S8460 = 8460;
  localparam test_b1_S8461 = 8461;
  localparam test_b1_S8462 = 8462;
  localparam test_b1_S8463 = 8463;
  localparam test_b1_S8464 = 8464;
  localparam test_b1_S8465 = 8465;
  localparam test_b1_S8466 = 8466;
  localparam test_b1_S8467 = 8467;
  localparam test_b1_S8468 = 8468;
  localparam test_b1_S8469 = 8469;
  localparam test_b1_S8470 = 8470;
  localparam test_b1_S8471 = 8471;
  localparam test_b1_S8472 = 8472;
  localparam test_b1_S8473 = 8473;
  localparam test_b1_S8474 = 8474;
  localparam test_b1_S8475 = 8475;
  localparam test_b1_S8476 = 8476;
  localparam test_b1_S8477 = 8477;
  localparam test_b1_S8478 = 8478;
  localparam test_b1_S8479 = 8479;
  localparam test_b1_S8480 = 8480;
  localparam test_b1_S8481 = 8481;
  localparam test_b1_S8482 = 8482;
  localparam test_b1_S8483 = 8483;
  localparam test_b1_S8484 = 8484;
  localparam test_b1_S8485 = 8485;
  localparam test_b1_S8486 = 8486;
  localparam test_b1_S8487 = 8487;
  localparam test_b1_S8488 = 8488;
  localparam test_b1_S8489 = 8489;
  localparam test_b1_S8490 = 8490;
  localparam test_b1_S8491 = 8491;
  localparam test_b1_S8492 = 8492;
  localparam test_b1_S8493 = 8493;
  localparam test_b1_S8494 = 8494;
  localparam test_b1_S8495 = 8495;
  localparam test_b1_S8496 = 8496;
  localparam test_b1_S8497 = 8497;
  localparam test_b1_S8498 = 8498;
  localparam test_b1_S8499 = 8499;
  localparam test_b1_S8500 = 8500;
  localparam test_b1_S8501 = 8501;
  localparam test_b1_S8502 = 8502;
  localparam test_b1_S8503 = 8503;
  localparam test_b1_S8504 = 8504;
  localparam test_b1_S8505 = 8505;
  localparam test_b1_S8506 = 8506;
  localparam test_b1_S8507 = 8507;
  localparam test_b1_S8508 = 8508;
  localparam test_b1_S8509 = 8509;
  localparam test_b1_S8510 = 8510;
  localparam test_b1_S8511 = 8511;
  localparam test_b1_S8512 = 8512;
  localparam test_b1_S8513 = 8513;
  localparam test_b1_S8514 = 8514;
  localparam test_b1_S8515 = 8515;
  localparam test_b1_S8516 = 8516;
  localparam test_b1_S8517 = 8517;
  localparam test_b1_S8518 = 8518;
  localparam test_b1_S8519 = 8519;
  localparam test_b1_S8520 = 8520;
  localparam test_b1_S8521 = 8521;
  localparam test_b1_S8522 = 8522;
  localparam test_b1_S8523 = 8523;
  localparam test_b1_S8524 = 8524;
  localparam test_b1_S8525 = 8525;
  localparam test_b1_S8526 = 8526;
  localparam test_b1_S8527 = 8527;
  localparam test_b1_S8528 = 8528;
  localparam test_b1_S8529 = 8529;
  localparam test_b1_S8530 = 8530;
  localparam test_b1_S8531 = 8531;
  localparam test_b1_S8532 = 8532;
  localparam test_b1_S8533 = 8533;
  localparam test_b1_S8534 = 8534;
  localparam test_b1_S8535 = 8535;
  localparam test_b1_S8536 = 8536;
  localparam test_b1_S8537 = 8537;
  localparam test_b1_S8538 = 8538;
  localparam test_b1_S8539 = 8539;
  localparam test_b1_S8540 = 8540;
  localparam test_b1_S8541 = 8541;
  localparam test_b1_S8542 = 8542;
  localparam test_b1_S8543 = 8543;
  localparam test_b1_S8544 = 8544;
  localparam test_b1_S8545 = 8545;
  localparam test_b1_S8546 = 8546;
  localparam test_b1_S8547 = 8547;
  localparam test_b1_S8548 = 8548;
  localparam test_b1_S8549 = 8549;
  localparam test_b1_S8550 = 8550;
  localparam test_b1_S8551 = 8551;
  localparam test_b1_S8552 = 8552;
  localparam test_b1_S8553 = 8553;
  localparam test_b1_FINISH = 8554;
  
  //signals: 
  wire retro_main_0_valid;
  reg clk;
  reg retro_main_0_accept;
  reg retro_main_0_ready;
  reg rst;
  reg        [13:0] test_state;
  //signals: IMAGE
  wire        [14:0] IMAGE_len;
  wire        [31:0] IMAGE_q;
  reg        [14:0] IMAGE_addr;
  reg        [31:0] IMAGE_d;
  reg IMAGE_req;
  reg IMAGE_we;
  //signals: in_io_ports
  wire        [4:0] retro_main_0_in_io_ports_addr;
  wire        [31:0] retro_main_0_in_io_ports_d;
  wire        [4:0] retro_main_0_in_io_ports_len;
  wire        [31:0] retro_main_0_in_io_ports_q;
  wire retro_main_0_in_io_ports_req;
  wire retro_main_0_in_io_ports_we;
  //signals: in_memory
  wire        [14:0] retro_main_0_in_memory_addr;
  wire        [31:0] retro_main_0_in_memory_d;
  wire        [14:0] retro_main_0_in_memory_len;
  wire        [31:0] retro_main_0_in_memory_q;
  wire retro_main_0_in_memory_req;
  wire retro_main_0_in_memory_we;
  //signals: io_ports
  wire        [4:0] io_ports_len;
  wire        [31:0] io_ports_q;
  reg        [4:0] io_ports_addr;
  reg        [31:0] io_ports_d;
  reg io_ports_req;
  reg io_ports_we;
  //signals: o2n_array10012854
  wire        [1:0] o2n_array10012854_switch;
  //signals: o2n_array10022855
  wire        [1:0] o2n_array10022855_switch;
  //signals: ram
  wire        [4:0] array1001_ram_addr;
  wire        [31:0] array1001_ram_d;
  wire        [4:0] array1001_ram_len;
  wire        [31:0] array1001_ram_q;
  wire array1001_ram_we;
  wire        [14:0] array1002_ram_addr;
  wire        [31:0] array1002_ram_d;
  wire        [14:0] array1002_ram_len;
  wire        [31:0] array1002_ram_q;
  wire array1002_ram_we;
  //combinations: o2n_array10012854
  assign retro_main_0_in_io_ports_q = 1'b1 == o2n_array10012854_switch[0] ? array1001_ram_q:32'd0;
  assign io_ports_q = 1'b1 == o2n_array10012854_switch[1] ? array1001_ram_q:32'd0;
  assign array1001_ram_addr = 1'b1 == o2n_array10012854_switch[0] ? retro_main_0_in_io_ports_addr:
                              1'b1 == o2n_array10012854_switch[1] ? io_ports_addr:5'd0;
  assign array1001_ram_d = 1'b1 == o2n_array10012854_switch[0] ? retro_main_0_in_io_ports_d:
                           1'b1 == o2n_array10012854_switch[1] ? io_ports_d:32'd0;
  assign array1001_ram_we = 1'b1 == o2n_array10012854_switch[0] ? retro_main_0_in_io_ports_we:
                            1'b1 == o2n_array10012854_switch[1] ? io_ports_we:1'd0;
  assign io_ports_len = array1001_ram_len;
  assign o2n_array10012854_switch = {io_ports_req, retro_main_0_in_io_ports_req};
  assign retro_main_0_in_io_ports_len = array1001_ram_len;
  //combinations: o2n_array10022855
  assign retro_main_0_in_memory_q = 1'b1 == o2n_array10022855_switch[0] ? array1002_ram_q:32'd0;
  assign IMAGE_q = 1'b1 == o2n_array10022855_switch[1] ? array1002_ram_q:32'd0;
  assign IMAGE_len = array1002_ram_len;
  assign array1002_ram_addr = 1'b1 == o2n_array10022855_switch[0] ? retro_main_0_in_memory_addr:
                              1'b1 == o2n_array10022855_switch[1] ? IMAGE_addr:15'd0;
  assign array1002_ram_d = 1'b1 == o2n_array10022855_switch[0] ? retro_main_0_in_memory_d:
                           1'b1 == o2n_array10022855_switch[1] ? IMAGE_d:32'd0;
  assign array1002_ram_we = 1'b1 == o2n_array10022855_switch[0] ? retro_main_0_in_memory_we:
                            1'b1 == o2n_array10022855_switch[1] ? IMAGE_we:1'd0;
  assign o2n_array10022855_switch = {IMAGE_req, retro_main_0_in_memory_req};
  assign retro_main_0_in_memory_len = array1002_ram_len;
  //sub modules
  //array1001 instance
  BidirectionalSinglePortRam#(
    .DATA_WIDTH(32),
    .ADDR_WIDTH(5),
    .RAM_LENGTH(16)
    )
    array1001(
      .clk(clk),
      .rst(rst),
      .ram_addr(array1001_ram_addr),
      .ram_d(array1001_ram_d),
      .ram_we(array1001_ram_we),
      .ram_q(array1001_ram_q),
      .ram_len(array1001_ram_len)
    );
  //array1002 instance
  BidirectionalSinglePortRam#(
    .DATA_WIDTH(32),
    .ADDR_WIDTH(15),
    .RAM_LENGTH(8533)
    )
    array1002(
      .clk(clk),
      .rst(rst),
      .ram_addr(array1002_ram_addr),
      .ram_d(array1002_ram_d),
      .ram_we(array1002_ram_we),
      .ram_q(array1002_ram_q),
      .ram_len(array1002_ram_len)
    );
  //retro_main_0 instance
  retro_main retro_main_0(
    .clk(clk),
    .rst(rst),
    .retro_main_ready(retro_main_0_ready),
    .retro_main_accept(retro_main_0_accept),
    .retro_main_valid(retro_main_0_valid),
    .retro_main_in_memory_addr(retro_main_0_in_memory_addr),
    .retro_main_in_memory_d(retro_main_0_in_memory_d),
    .retro_main_in_memory_we(retro_main_0_in_memory_we),
    .retro_main_in_memory_q(retro_main_0_in_memory_q),
    .retro_main_in_memory_len(retro_main_0_in_memory_len),
    .retro_main_in_memory_req(retro_main_0_in_memory_req),
    .retro_main_in_io_ports_addr(retro_main_0_in_io_ports_addr),
    .retro_main_in_io_ports_d(retro_main_0_in_io_ports_d),
    .retro_main_in_io_ports_we(retro_main_0_in_io_ports_we),
    .retro_main_in_io_ports_q(retro_main_0_in_io_ports_q),
    .retro_main_in_io_ports_len(retro_main_0_in_io_ports_len),
    .retro_main_in_io_ports_req(retro_main_0_in_io_ports_req)
  );
  
  
  initial begin
    clk = 0;
    #CLK_HALF_PERIOD
    forever #CLK_HALF_PERIOD clk = ~clk;
  end
  initial begin
    rst <= 1;
    #INITIAL_RESET_SPAN
    rst <= 0;
  end
  

  always @(posedge clk) begin
    if (rst) begin
      IMAGE_addr <= 0;
      IMAGE_d <= 0;
      IMAGE_req <= 0;
      IMAGE_we <= 0;
      io_ports_addr <= 0;
      io_ports_d <= 0;
      io_ports_req <= 0;
      io_ports_we <= 0;
      retro_main_0_accept <= 0;
      retro_main_0_ready <= 0;
      test_state <= test_b1_INIT;
    end else begin //if (rst)
      case(test_state)
      test_b1_INIT: begin
        io_ports_addr <= 0;
        io_ports_we <= 1;
        io_ports_req <= 1;
        io_ports_d <= 0;
        test_state <= test_b1_S1;
      end
      test_b1_S1: begin
        io_ports_addr <= 1;
        io_ports_we <= 1;
        io_ports_req <= 1;
        io_ports_d <= 0;
        test_state <= test_b1_S2;
      end
      test_b1_S2: begin
        io_ports_addr <= 2;
        io_ports_we <= 1;
        io_ports_req <= 1;
        io_ports_d <= 0;
        test_state <= test_b1_S3;
      end
      test_b1_S3: begin
        io_ports_addr <= 3;
        io_ports_we <= 1;
        io_ports_req <= 1;
        io_ports_d <= 0;
        test_state <= test_b1_S4;
      end
      test_b1_S4: begin
        io_ports_addr <= 4;
        io_ports_we <= 1;
        io_ports_req <= 1;
        io_ports_d <= 0;
        test_state <= test_b1_S5;
      end
      test_b1_S5: begin
        io_ports_addr <= 5;
        io_ports_we <= 1;
        io_ports_req <= 1;
        io_ports_d <= 0;
        test_state <= test_b1_S6;
      end
      test_b1_S6: begin
        io_ports_addr <= 6;
        io_ports_we <= 1;
        io_ports_req <= 1;
        io_ports_d <= 0;
        test_state <= test_b1_S7;
      end
      test_b1_S7: begin
        io_ports_addr <= 7;
        io_ports_we <= 1;
        io_ports_req <= 1;
        io_ports_d <= 0;
        test_state <= test_b1_S8;
      end
      test_b1_S8: begin
        io_ports_addr <= 8;
        io_ports_we <= 1;
        io_ports_req <= 1;
        io_ports_d <= 0;
        test_state <= test_b1_S9;
      end
      test_b1_S9: begin
        io_ports_addr <= 9;
        io_ports_we <= 1;
        io_ports_req <= 1;
        io_ports_d <= 0;
        test_state <= test_b1_S10;
      end
      test_b1_S10: begin
        io_ports_addr <= 10;
        io_ports_we <= 1;
        io_ports_req <= 1;
        io_ports_d <= 0;
        test_state <= test_b1_S11;
      end
      test_b1_S11: begin
        io_ports_addr <= 11;
        io_ports_we <= 1;
        io_ports_req <= 1;
        io_ports_d <= 0;
        test_state <= test_b1_S12;
      end
      test_b1_S12: begin
        io_ports_addr <= 12;
        io_ports_we <= 1;
        io_ports_req <= 1;
        io_ports_d <= 0;
        test_state <= test_b1_S13;
      end
      test_b1_S13: begin
        io_ports_addr <= 13;
        io_ports_we <= 1;
        io_ports_req <= 1;
        io_ports_d <= 0;
        test_state <= test_b1_S14;
      end
      test_b1_S14: begin
        io_ports_addr <= 14;
        io_ports_we <= 1;
        io_ports_req <= 1;
        io_ports_d <= 0;
        test_state <= test_b1_S15;
      end
      test_b1_S15: begin
        io_ports_addr <= 15;
        io_ports_we <= 1;
        io_ports_req <= 1;
        io_ports_d <= 0;
        test_state <= test_b1_S16;
      end
      test_b1_S16: begin
        IMAGE_addr <= 0;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8;
        io_ports_req <= 0;
        test_state <= test_b1_S17;
      end
      test_b1_S17: begin
        IMAGE_addr <= 1;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2311;
        test_state <= test_b1_S18;
      end
      test_b1_S18: begin
        IMAGE_addr <= 2;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8479;
        test_state <= test_b1_S19;
      end
      test_b1_S19: begin
        IMAGE_addr <= 3;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8533;
        test_state <= test_b1_S20;
      end
      test_b1_S20: begin
        IMAGE_addr <= 4;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S21;
      end
      test_b1_S21: begin
        IMAGE_addr <= 5;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6503;
        test_state <= test_b1_S22;
      end
      test_b1_S22: begin
        IMAGE_addr <= 6;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2314;
        test_state <= test_b1_S23;
      end
      test_b1_S23: begin
        IMAGE_addr <= 7;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 82;
        test_state <= test_b1_S24;
      end
      test_b1_S24: begin
        IMAGE_addr <= 8;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S25;
      end
      test_b1_S25: begin
        IMAGE_addr <= 9;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S26;
      end
      test_b1_S26: begin
        IMAGE_addr <= 10;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S27;
      end
      test_b1_S27: begin
        IMAGE_addr <= 11;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 111;
        test_state <= test_b1_S28;
      end
      test_b1_S28: begin
        IMAGE_addr <= 12;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S29;
      end
      test_b1_S29: begin
        IMAGE_addr <= 13;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 49;
        test_state <= test_b1_S30;
      end
      test_b1_S30: begin
        IMAGE_addr <= 14;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 49;
        test_state <= test_b1_S31;
      end
      test_b1_S31: begin
        IMAGE_addr <= 15;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 46;
        test_state <= test_b1_S32;
      end
      test_b1_S32: begin
        IMAGE_addr <= 16;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 52;
        test_state <= test_b1_S33;
      end
      test_b1_S33: begin
        IMAGE_addr <= 17;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S34;
      end
      test_b1_S34: begin
        IMAGE_addr <= 18;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 50;
        test_state <= test_b1_S35;
      end
      test_b1_S35: begin
        IMAGE_addr <= 19;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 48;
        test_state <= test_b1_S36;
      end
      test_b1_S36: begin
        IMAGE_addr <= 20;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 49;
        test_state <= test_b1_S37;
      end
      test_b1_S37: begin
        IMAGE_addr <= 21;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 50;
        test_state <= test_b1_S38;
      end
      test_b1_S38: begin
        IMAGE_addr <= 22;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 46;
        test_state <= test_b1_S39;
      end
      test_b1_S39: begin
        IMAGE_addr <= 23;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 48;
        test_state <= test_b1_S40;
      end
      test_b1_S40: begin
        IMAGE_addr <= 24;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 51;
        test_state <= test_b1_S41;
      end
      test_b1_S41: begin
        IMAGE_addr <= 25;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 46;
        test_state <= test_b1_S42;
      end
      test_b1_S42: begin
        IMAGE_addr <= 26;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 49;
        test_state <= test_b1_S43;
      end
      test_b1_S43: begin
        IMAGE_addr <= 27;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 57;
        test_state <= test_b1_S44;
      end
      test_b1_S44: begin
        IMAGE_addr <= 28;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S45;
      end
      test_b1_S45: begin
        IMAGE_addr <= 29;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 111;
        test_state <= test_b1_S46;
      end
      test_b1_S46: begin
        IMAGE_addr <= 30;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 107;
        test_state <= test_b1_S47;
      end
      test_b1_S47: begin
        IMAGE_addr <= 31;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 32;
        test_state <= test_b1_S48;
      end
      test_b1_S48: begin
        IMAGE_addr <= 32;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S49;
      end
      test_b1_S49: begin
        IMAGE_addr <= 33;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S50;
      end
      test_b1_S50: begin
        IMAGE_addr <= 34;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S51;
      end
      test_b1_S51: begin
        IMAGE_addr <= 35;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S52;
      end
      test_b1_S52: begin
        IMAGE_addr <= 36;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S53;
      end
      test_b1_S53: begin
        IMAGE_addr <= 37;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S54;
      end
      test_b1_S54: begin
        IMAGE_addr <= 38;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S55;
      end
      test_b1_S55: begin
        IMAGE_addr <= 39;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 26;
        test_state <= test_b1_S56;
      end
      test_b1_S56: begin
        IMAGE_addr <= 40;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S57;
      end
      test_b1_S57: begin
        IMAGE_addr <= 41;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S58;
      end
      test_b1_S58: begin
        IMAGE_addr <= 42;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S59;
      end
      test_b1_S59: begin
        IMAGE_addr <= 43;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S60;
      end
      test_b1_S60: begin
        IMAGE_addr <= 44;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 27;
        test_state <= test_b1_S61;
      end
      test_b1_S61: begin
        IMAGE_addr <= 45;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S62;
      end
      test_b1_S62: begin
        IMAGE_addr <= 46;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S63;
      end
      test_b1_S63: begin
        IMAGE_addr <= 47;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S64;
      end
      test_b1_S64: begin
        IMAGE_addr <= 48;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S65;
      end
      test_b1_S65: begin
        IMAGE_addr <= 49;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S66;
      end
      test_b1_S66: begin
        IMAGE_addr <= 50;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S67;
      end
      test_b1_S67: begin
        IMAGE_addr <= 51;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S68;
      end
      test_b1_S68: begin
        IMAGE_addr <= 52;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S69;
      end
      test_b1_S69: begin
        IMAGE_addr <= 53;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S70;
      end
      test_b1_S70: begin
        IMAGE_addr <= 54;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S71;
      end
      test_b1_S71: begin
        IMAGE_addr <= 55;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S72;
      end
      test_b1_S72: begin
        IMAGE_addr <= 56;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S73;
      end
      test_b1_S73: begin
        IMAGE_addr <= 57;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S74;
      end
      test_b1_S74: begin
        IMAGE_addr <= 58;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S75;
      end
      test_b1_S75: begin
        IMAGE_addr <= 59;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 20;
        test_state <= test_b1_S76;
      end
      test_b1_S76: begin
        IMAGE_addr <= 60;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S77;
      end
      test_b1_S77: begin
        IMAGE_addr <= 61;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S78;
      end
      test_b1_S78: begin
        IMAGE_addr <= 62;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S79;
      end
      test_b1_S79: begin
        IMAGE_addr <= 63;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S80;
      end
      test_b1_S80: begin
        IMAGE_addr <= 64;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 21;
        test_state <= test_b1_S81;
      end
      test_b1_S81: begin
        IMAGE_addr <= 65;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S82;
      end
      test_b1_S82: begin
        IMAGE_addr <= 66;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S83;
      end
      test_b1_S83: begin
        IMAGE_addr <= 67;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S84;
      end
      test_b1_S84: begin
        IMAGE_addr <= 68;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S85;
      end
      test_b1_S85: begin
        IMAGE_addr <= 69;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 22;
        test_state <= test_b1_S86;
      end
      test_b1_S86: begin
        IMAGE_addr <= 70;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S87;
      end
      test_b1_S87: begin
        IMAGE_addr <= 71;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S88;
      end
      test_b1_S88: begin
        IMAGE_addr <= 72;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S89;
      end
      test_b1_S89: begin
        IMAGE_addr <= 73;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S90;
      end
      test_b1_S90: begin
        IMAGE_addr <= 74;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S91;
      end
      test_b1_S91: begin
        IMAGE_addr <= 75;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S92;
      end
      test_b1_S92: begin
        IMAGE_addr <= 76;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S93;
      end
      test_b1_S93: begin
        IMAGE_addr <= 77;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S94;
      end
      test_b1_S94: begin
        IMAGE_addr <= 78;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S95;
      end
      test_b1_S95: begin
        IMAGE_addr <= 79;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S96;
      end
      test_b1_S96: begin
        IMAGE_addr <= 80;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S97;
      end
      test_b1_S97: begin
        IMAGE_addr <= 81;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S98;
      end
      test_b1_S98: begin
        IMAGE_addr <= 82;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S99;
      end
      test_b1_S99: begin
        IMAGE_addr <= 83;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S100;
      end
      test_b1_S100: begin
        IMAGE_addr <= 84;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 16;
        test_state <= test_b1_S101;
      end
      test_b1_S101: begin
        IMAGE_addr <= 85;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S102;
      end
      test_b1_S102: begin
        IMAGE_addr <= 86;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S103;
      end
      test_b1_S103: begin
        IMAGE_addr <= 87;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S104;
      end
      test_b1_S104: begin
        IMAGE_addr <= 88;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S105;
      end
      test_b1_S105: begin
        IMAGE_addr <= 89;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 17;
        test_state <= test_b1_S106;
      end
      test_b1_S106: begin
        IMAGE_addr <= 90;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S107;
      end
      test_b1_S107: begin
        IMAGE_addr <= 91;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S108;
      end
      test_b1_S108: begin
        IMAGE_addr <= 92;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S109;
      end
      test_b1_S109: begin
        IMAGE_addr <= 93;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S110;
      end
      test_b1_S110: begin
        IMAGE_addr <= 94;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 18;
        test_state <= test_b1_S111;
      end
      test_b1_S111: begin
        IMAGE_addr <= 95;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S112;
      end
      test_b1_S112: begin
        IMAGE_addr <= 96;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S113;
      end
      test_b1_S113: begin
        IMAGE_addr <= 97;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S114;
      end
      test_b1_S114: begin
        IMAGE_addr <= 98;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S115;
      end
      test_b1_S115: begin
        IMAGE_addr <= 99;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 19;
        test_state <= test_b1_S116;
      end
      test_b1_S116: begin
        IMAGE_addr <= 100;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S117;
      end
      test_b1_S117: begin
        IMAGE_addr <= 101;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S118;
      end
      test_b1_S118: begin
        IMAGE_addr <= 102;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S119;
      end
      test_b1_S119: begin
        IMAGE_addr <= 103;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S120;
      end
      test_b1_S120: begin
        IMAGE_addr <= 104;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 23;
        test_state <= test_b1_S121;
      end
      test_b1_S121: begin
        IMAGE_addr <= 105;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S122;
      end
      test_b1_S122: begin
        IMAGE_addr <= 106;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S123;
      end
      test_b1_S123: begin
        IMAGE_addr <= 107;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S124;
      end
      test_b1_S124: begin
        IMAGE_addr <= 108;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S125;
      end
      test_b1_S125: begin
        IMAGE_addr <= 109;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 24;
        test_state <= test_b1_S126;
      end
      test_b1_S126: begin
        IMAGE_addr <= 110;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S127;
      end
      test_b1_S127: begin
        IMAGE_addr <= 111;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S128;
      end
      test_b1_S128: begin
        IMAGE_addr <= 112;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S129;
      end
      test_b1_S129: begin
        IMAGE_addr <= 113;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S130;
      end
      test_b1_S130: begin
        IMAGE_addr <= 114;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 29;
        test_state <= test_b1_S131;
      end
      test_b1_S131: begin
        IMAGE_addr <= 115;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S132;
      end
      test_b1_S132: begin
        IMAGE_addr <= 116;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S133;
      end
      test_b1_S133: begin
        IMAGE_addr <= 117;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S134;
      end
      test_b1_S134: begin
        IMAGE_addr <= 118;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S135;
      end
      test_b1_S135: begin
        IMAGE_addr <= 119;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 28;
        test_state <= test_b1_S136;
      end
      test_b1_S136: begin
        IMAGE_addr <= 120;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S137;
      end
      test_b1_S137: begin
        IMAGE_addr <= 121;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S138;
      end
      test_b1_S138: begin
        IMAGE_addr <= 122;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S139;
      end
      test_b1_S139: begin
        IMAGE_addr <= 123;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S140;
      end
      test_b1_S140: begin
        IMAGE_addr <= 124;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S141;
      end
      test_b1_S141: begin
        IMAGE_addr <= 125;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S142;
      end
      test_b1_S142: begin
        IMAGE_addr <= 126;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S143;
      end
      test_b1_S143: begin
        IMAGE_addr <= 127;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S144;
      end
      test_b1_S144: begin
        IMAGE_addr <= 128;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 29;
        test_state <= test_b1_S145;
      end
      test_b1_S145: begin
        IMAGE_addr <= 129;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 30;
        test_state <= test_b1_S146;
      end
      test_b1_S146: begin
        IMAGE_addr <= 130;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S147;
      end
      test_b1_S147: begin
        IMAGE_addr <= 131;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S148;
      end
      test_b1_S148: begin
        IMAGE_addr <= 132;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S149;
      end
      test_b1_S149: begin
        IMAGE_addr <= 133;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S150;
      end
      test_b1_S150: begin
        IMAGE_addr <= 134;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5;
        test_state <= test_b1_S151;
      end
      test_b1_S151: begin
        IMAGE_addr <= 135;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S152;
      end
      test_b1_S152: begin
        IMAGE_addr <= 136;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6;
        test_state <= test_b1_S153;
      end
      test_b1_S153: begin
        IMAGE_addr <= 137;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S154;
      end
      test_b1_S154: begin
        IMAGE_addr <= 138;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S155;
      end
      test_b1_S155: begin
        IMAGE_addr <= 139;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S156;
      end
      test_b1_S156: begin
        IMAGE_addr <= 140;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S157;
      end
      test_b1_S157: begin
        IMAGE_addr <= 141;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S158;
      end
      test_b1_S158: begin
        IMAGE_addr <= 142;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S159;
      end
      test_b1_S159: begin
        IMAGE_addr <= 143;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4294967295;
        test_state <= test_b1_S160;
      end
      test_b1_S160: begin
        IMAGE_addr <= 144;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 22;
        test_state <= test_b1_S161;
      end
      test_b1_S161: begin
        IMAGE_addr <= 145;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S162;
      end
      test_b1_S162: begin
        IMAGE_addr <= 146;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S163;
      end
      test_b1_S163: begin
        IMAGE_addr <= 147;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S164;
      end
      test_b1_S164: begin
        IMAGE_addr <= 148;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S165;
      end
      test_b1_S165: begin
        IMAGE_addr <= 149;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S166;
      end
      test_b1_S166: begin
        IMAGE_addr <= 150;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4294967295;
        test_state <= test_b1_S167;
      end
      test_b1_S167: begin
        IMAGE_addr <= 151;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S168;
      end
      test_b1_S168: begin
        IMAGE_addr <= 152;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S169;
      end
      test_b1_S169: begin
        IMAGE_addr <= 153;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S170;
      end
      test_b1_S170: begin
        IMAGE_addr <= 154;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S171;
      end
      test_b1_S171: begin
        IMAGE_addr <= 155;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S172;
      end
      test_b1_S172: begin
        IMAGE_addr <= 156;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S173;
      end
      test_b1_S173: begin
        IMAGE_addr <= 157;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S174;
      end
      test_b1_S174: begin
        IMAGE_addr <= 158;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S175;
      end
      test_b1_S175: begin
        IMAGE_addr <= 159;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S176;
      end
      test_b1_S176: begin
        IMAGE_addr <= 160;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S177;
      end
      test_b1_S177: begin
        IMAGE_addr <= 161;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S178;
      end
      test_b1_S178: begin
        IMAGE_addr <= 162;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S179;
      end
      test_b1_S179: begin
        IMAGE_addr <= 163;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S180;
      end
      test_b1_S180: begin
        IMAGE_addr <= 164;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S181;
      end
      test_b1_S181: begin
        IMAGE_addr <= 165;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 19;
        test_state <= test_b1_S182;
      end
      test_b1_S182: begin
        IMAGE_addr <= 166;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S183;
      end
      test_b1_S183: begin
        IMAGE_addr <= 167;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S184;
      end
      test_b1_S184: begin
        IMAGE_addr <= 168;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S185;
      end
      test_b1_S185: begin
        IMAGE_addr <= 169;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S186;
      end
      test_b1_S186: begin
        IMAGE_addr <= 170;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S187;
      end
      test_b1_S187: begin
        IMAGE_addr <= 171;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S188;
      end
      test_b1_S188: begin
        IMAGE_addr <= 172;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 19;
        test_state <= test_b1_S189;
      end
      test_b1_S189: begin
        IMAGE_addr <= 173;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S190;
      end
      test_b1_S190: begin
        IMAGE_addr <= 174;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S191;
      end
      test_b1_S191: begin
        IMAGE_addr <= 175;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S192;
      end
      test_b1_S192: begin
        IMAGE_addr <= 176;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S193;
      end
      test_b1_S193: begin
        IMAGE_addr <= 177;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S194;
      end
      test_b1_S194: begin
        IMAGE_addr <= 178;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S195;
      end
      test_b1_S195: begin
        IMAGE_addr <= 179;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4294967295;
        test_state <= test_b1_S196;
      end
      test_b1_S196: begin
        IMAGE_addr <= 180;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 18;
        test_state <= test_b1_S197;
      end
      test_b1_S197: begin
        IMAGE_addr <= 181;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S198;
      end
      test_b1_S198: begin
        IMAGE_addr <= 182;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S199;
      end
      test_b1_S199: begin
        IMAGE_addr <= 183;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S200;
      end
      test_b1_S200: begin
        IMAGE_addr <= 184;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S201;
      end
      test_b1_S201: begin
        IMAGE_addr <= 185;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 27;
        test_state <= test_b1_S202;
      end
      test_b1_S202: begin
        IMAGE_addr <= 186;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5;
        test_state <= test_b1_S203;
      end
      test_b1_S203: begin
        IMAGE_addr <= 187;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S204;
      end
      test_b1_S204: begin
        IMAGE_addr <= 188;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S205;
      end
      test_b1_S205: begin
        IMAGE_addr <= 189;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S206;
      end
      test_b1_S206: begin
        IMAGE_addr <= 190;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S207;
      end
      test_b1_S207: begin
        IMAGE_addr <= 191;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S208;
      end
      test_b1_S208: begin
        IMAGE_addr <= 192;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 26;
        test_state <= test_b1_S209;
      end
      test_b1_S209: begin
        IMAGE_addr <= 193;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S210;
      end
      test_b1_S210: begin
        IMAGE_addr <= 194;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S211;
      end
      test_b1_S211: begin
        IMAGE_addr <= 195;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S212;
      end
      test_b1_S212: begin
        IMAGE_addr <= 196;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S213;
      end
      test_b1_S213: begin
        IMAGE_addr <= 197;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S214;
      end
      test_b1_S214: begin
        IMAGE_addr <= 198;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S215;
      end
      test_b1_S215: begin
        IMAGE_addr <= 199;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S216;
      end
      test_b1_S216: begin
        IMAGE_addr <= 200;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 26;
        test_state <= test_b1_S217;
      end
      test_b1_S217: begin
        IMAGE_addr <= 201;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5;
        test_state <= test_b1_S218;
      end
      test_b1_S218: begin
        IMAGE_addr <= 202;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S219;
      end
      test_b1_S219: begin
        IMAGE_addr <= 203;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6;
        test_state <= test_b1_S220;
      end
      test_b1_S220: begin
        IMAGE_addr <= 204;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S221;
      end
      test_b1_S221: begin
        IMAGE_addr <= 205;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S222;
      end
      test_b1_S222: begin
        IMAGE_addr <= 206;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S223;
      end
      test_b1_S223: begin
        IMAGE_addr <= 207;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S224;
      end
      test_b1_S224: begin
        IMAGE_addr <= 208;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S225;
      end
      test_b1_S225: begin
        IMAGE_addr <= 209;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S226;
      end
      test_b1_S226: begin
        IMAGE_addr <= 210;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S227;
      end
      test_b1_S227: begin
        IMAGE_addr <= 211;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S228;
      end
      test_b1_S228: begin
        IMAGE_addr <= 212;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S229;
      end
      test_b1_S229: begin
        IMAGE_addr <= 213;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S230;
      end
      test_b1_S230: begin
        IMAGE_addr <= 214;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S231;
      end
      test_b1_S231: begin
        IMAGE_addr <= 215;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 206;
        test_state <= test_b1_S232;
      end
      test_b1_S232: begin
        IMAGE_addr <= 216;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 197;
        test_state <= test_b1_S233;
      end
      test_b1_S233: begin
        IMAGE_addr <= 217;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S234;
      end
      test_b1_S234: begin
        IMAGE_addr <= 218;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S235;
      end
      test_b1_S235: begin
        IMAGE_addr <= 219;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S236;
      end
      test_b1_S236: begin
        IMAGE_addr <= 220;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S237;
      end
      test_b1_S237: begin
        IMAGE_addr <= 221;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S238;
      end
      test_b1_S238: begin
        IMAGE_addr <= 222;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S239;
      end
      test_b1_S239: begin
        IMAGE_addr <= 223;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S240;
      end
      test_b1_S240: begin
        IMAGE_addr <= 224;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S241;
      end
      test_b1_S241: begin
        IMAGE_addr <= 225;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S242;
      end
      test_b1_S242: begin
        IMAGE_addr <= 226;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 213;
        test_state <= test_b1_S243;
      end
      test_b1_S243: begin
        IMAGE_addr <= 227;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S244;
      end
      test_b1_S244: begin
        IMAGE_addr <= 228;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S245;
      end
      test_b1_S245: begin
        IMAGE_addr <= 229;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S246;
      end
      test_b1_S246: begin
        IMAGE_addr <= 230;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S247;
      end
      test_b1_S247: begin
        IMAGE_addr <= 231;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 222;
        test_state <= test_b1_S248;
      end
      test_b1_S248: begin
        IMAGE_addr <= 232;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 222;
        test_state <= test_b1_S249;
      end
      test_b1_S249: begin
        IMAGE_addr <= 233;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S250;
      end
      test_b1_S250: begin
        IMAGE_addr <= 234;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S251;
      end
      test_b1_S251: begin
        IMAGE_addr <= 235;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 155;
        test_state <= test_b1_S252;
      end
      test_b1_S252: begin
        IMAGE_addr <= 236;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S253;
      end
      test_b1_S253: begin
        IMAGE_addr <= 237;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S254;
      end
      test_b1_S254: begin
        IMAGE_addr <= 238;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 189;
        test_state <= test_b1_S255;
      end
      test_b1_S255: begin
        IMAGE_addr <= 239;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 25;
        test_state <= test_b1_S256;
      end
      test_b1_S256: begin
        IMAGE_addr <= 240;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 213;
        test_state <= test_b1_S257;
      end
      test_b1_S257: begin
        IMAGE_addr <= 241;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8;
        test_state <= test_b1_S258;
      end
      test_b1_S258: begin
        IMAGE_addr <= 242;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 238;
        test_state <= test_b1_S259;
      end
      test_b1_S259: begin
        IMAGE_addr <= 243;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S260;
      end
      test_b1_S260: begin
        IMAGE_addr <= 244;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S261;
      end
      test_b1_S261: begin
        IMAGE_addr <= 245;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 238;
        test_state <= test_b1_S262;
      end
      test_b1_S262: begin
        IMAGE_addr <= 246;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S263;
      end
      test_b1_S263: begin
        IMAGE_addr <= 247;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S264;
      end
      test_b1_S264: begin
        IMAGE_addr <= 248;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S265;
      end
      test_b1_S265: begin
        IMAGE_addr <= 249;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 213;
        test_state <= test_b1_S266;
      end
      test_b1_S266: begin
        IMAGE_addr <= 250;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S267;
      end
      test_b1_S267: begin
        IMAGE_addr <= 251;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S268;
      end
      test_b1_S268: begin
        IMAGE_addr <= 252;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S269;
      end
      test_b1_S269: begin
        IMAGE_addr <= 253;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S270;
      end
      test_b1_S270: begin
        IMAGE_addr <= 254;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S271;
      end
      test_b1_S271: begin
        IMAGE_addr <= 255;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5;
        test_state <= test_b1_S272;
      end
      test_b1_S272: begin
        IMAGE_addr <= 256;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 213;
        test_state <= test_b1_S273;
      end
      test_b1_S273: begin
        IMAGE_addr <= 257;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S274;
      end
      test_b1_S274: begin
        IMAGE_addr <= 258;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S275;
      end
      test_b1_S275: begin
        IMAGE_addr <= 259;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S276;
      end
      test_b1_S276: begin
        IMAGE_addr <= 260;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S277;
      end
      test_b1_S277: begin
        IMAGE_addr <= 261;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S278;
      end
      test_b1_S278: begin
        IMAGE_addr <= 262;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6;
        test_state <= test_b1_S279;
      end
      test_b1_S279: begin
        IMAGE_addr <= 263;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 213;
        test_state <= test_b1_S280;
      end
      test_b1_S280: begin
        IMAGE_addr <= 264;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S281;
      end
      test_b1_S281: begin
        IMAGE_addr <= 265;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S282;
      end
      test_b1_S282: begin
        IMAGE_addr <= 266;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S283;
      end
      test_b1_S283: begin
        IMAGE_addr <= 267;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S284;
      end
      test_b1_S284: begin
        IMAGE_addr <= 268;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S285;
      end
      test_b1_S285: begin
        IMAGE_addr <= 269;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 25;
        test_state <= test_b1_S286;
      end
      test_b1_S286: begin
        IMAGE_addr <= 270;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 213;
        test_state <= test_b1_S287;
      end
      test_b1_S287: begin
        IMAGE_addr <= 271;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S288;
      end
      test_b1_S288: begin
        IMAGE_addr <= 272;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S289;
      end
      test_b1_S289: begin
        IMAGE_addr <= 273;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S290;
      end
      test_b1_S290: begin
        IMAGE_addr <= 274;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S291;
      end
      test_b1_S291: begin
        IMAGE_addr <= 275;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 206;
        test_state <= test_b1_S292;
      end
      test_b1_S292: begin
        IMAGE_addr <= 276;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S293;
      end
      test_b1_S293: begin
        IMAGE_addr <= 277;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S294;
      end
      test_b1_S294: begin
        IMAGE_addr <= 278;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S295;
      end
      test_b1_S295: begin
        IMAGE_addr <= 279;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S296;
      end
      test_b1_S296: begin
        IMAGE_addr <= 280;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S297;
      end
      test_b1_S297: begin
        IMAGE_addr <= 281;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8;
        test_state <= test_b1_S298;
      end
      test_b1_S298: begin
        IMAGE_addr <= 282;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 213;
        test_state <= test_b1_S299;
      end
      test_b1_S299: begin
        IMAGE_addr <= 283;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 213;
        test_state <= test_b1_S300;
      end
      test_b1_S300: begin
        IMAGE_addr <= 284;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S301;
      end
      test_b1_S301: begin
        IMAGE_addr <= 285;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S302;
      end
      test_b1_S302: begin
        IMAGE_addr <= 286;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S303;
      end
      test_b1_S303: begin
        IMAGE_addr <= 287;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S304;
      end
      test_b1_S304: begin
        IMAGE_addr <= 288;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 27;
        test_state <= test_b1_S305;
      end
      test_b1_S305: begin
        IMAGE_addr <= 289;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5;
        test_state <= test_b1_S306;
      end
      test_b1_S306: begin
        IMAGE_addr <= 290;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S307;
      end
      test_b1_S307: begin
        IMAGE_addr <= 291;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S308;
      end
      test_b1_S308: begin
        IMAGE_addr <= 292;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S309;
      end
      test_b1_S309: begin
        IMAGE_addr <= 293;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S310;
      end
      test_b1_S310: begin
        IMAGE_addr <= 294;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S311;
      end
      test_b1_S311: begin
        IMAGE_addr <= 295;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S312;
      end
      test_b1_S312: begin
        IMAGE_addr <= 296;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S313;
      end
      test_b1_S313: begin
        IMAGE_addr <= 297;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S314;
      end
      test_b1_S314: begin
        IMAGE_addr <= 298;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S315;
      end
      test_b1_S315: begin
        IMAGE_addr <= 299;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 13;
        test_state <= test_b1_S316;
      end
      test_b1_S316: begin
        IMAGE_addr <= 300;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 304;
        test_state <= test_b1_S317;
      end
      test_b1_S317: begin
        IMAGE_addr <= 301;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 213;
        test_state <= test_b1_S318;
      end
      test_b1_S318: begin
        IMAGE_addr <= 302;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S319;
      end
      test_b1_S319: begin
        IMAGE_addr <= 303;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S320;
      end
      test_b1_S320: begin
        IMAGE_addr <= 304;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8;
        test_state <= test_b1_S321;
      end
      test_b1_S321: begin
        IMAGE_addr <= 305;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 183;
        test_state <= test_b1_S322;
      end
      test_b1_S322: begin
        IMAGE_addr <= 306;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S323;
      end
      test_b1_S323: begin
        IMAGE_addr <= 307;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S324;
      end
      test_b1_S324: begin
        IMAGE_addr <= 308;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8;
        test_state <= test_b1_S325;
      end
      test_b1_S325: begin
        IMAGE_addr <= 309;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 183;
        test_state <= test_b1_S326;
      end
      test_b1_S326: begin
        IMAGE_addr <= 310;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S327;
      end
      test_b1_S327: begin
        IMAGE_addr <= 311;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S328;
      end
      test_b1_S328: begin
        IMAGE_addr <= 312;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S329;
      end
      test_b1_S329: begin
        IMAGE_addr <= 313;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S330;
      end
      test_b1_S330: begin
        IMAGE_addr <= 314;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S331;
      end
      test_b1_S331: begin
        IMAGE_addr <= 315;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 25;
        test_state <= test_b1_S332;
      end
      test_b1_S332: begin
        IMAGE_addr <= 316;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S333;
      end
      test_b1_S333: begin
        IMAGE_addr <= 317;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S334;
      end
      test_b1_S334: begin
        IMAGE_addr <= 318;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S335;
      end
      test_b1_S335: begin
        IMAGE_addr <= 319;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 213;
        test_state <= test_b1_S336;
      end
      test_b1_S336: begin
        IMAGE_addr <= 320;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 213;
        test_state <= test_b1_S337;
      end
      test_b1_S337: begin
        IMAGE_addr <= 321;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S338;
      end
      test_b1_S338: begin
        IMAGE_addr <= 322;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S339;
      end
      test_b1_S339: begin
        IMAGE_addr <= 323;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S340;
      end
      test_b1_S340: begin
        IMAGE_addr <= 324;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S341;
      end
      test_b1_S341: begin
        IMAGE_addr <= 325;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S342;
      end
      test_b1_S342: begin
        IMAGE_addr <= 326;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S343;
      end
      test_b1_S343: begin
        IMAGE_addr <= 327;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S344;
      end
      test_b1_S344: begin
        IMAGE_addr <= 328;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S345;
      end
      test_b1_S345: begin
        IMAGE_addr <= 329;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 12;
        test_state <= test_b1_S346;
      end
      test_b1_S346: begin
        IMAGE_addr <= 330;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 342;
        test_state <= test_b1_S347;
      end
      test_b1_S347: begin
        IMAGE_addr <= 331;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S348;
      end
      test_b1_S348: begin
        IMAGE_addr <= 332;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S349;
      end
      test_b1_S349: begin
        IMAGE_addr <= 333;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S350;
      end
      test_b1_S350: begin
        IMAGE_addr <= 334;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S351;
      end
      test_b1_S351: begin
        IMAGE_addr <= 335;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4294967295;
        test_state <= test_b1_S352;
      end
      test_b1_S352: begin
        IMAGE_addr <= 336;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 12;
        test_state <= test_b1_S353;
      end
      test_b1_S353: begin
        IMAGE_addr <= 337;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 342;
        test_state <= test_b1_S354;
      end
      test_b1_S354: begin
        IMAGE_addr <= 338;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S355;
      end
      test_b1_S355: begin
        IMAGE_addr <= 339;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S356;
      end
      test_b1_S356: begin
        IMAGE_addr <= 340;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 16;
        test_state <= test_b1_S357;
      end
      test_b1_S357: begin
        IMAGE_addr <= 341;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S358;
      end
      test_b1_S358: begin
        IMAGE_addr <= 342;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8;
        test_state <= test_b1_S359;
      end
      test_b1_S359: begin
        IMAGE_addr <= 343;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S360;
      end
      test_b1_S360: begin
        IMAGE_addr <= 344;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4294967295;
        test_state <= test_b1_S361;
      end
      test_b1_S361: begin
        IMAGE_addr <= 345;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S362;
      end
      test_b1_S362: begin
        IMAGE_addr <= 346;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S363;
      end
      test_b1_S363: begin
        IMAGE_addr <= 347;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S364;
      end
      test_b1_S364: begin
        IMAGE_addr <= 348;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 344;
        test_state <= test_b1_S365;
      end
      test_b1_S365: begin
        IMAGE_addr <= 349;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S366;
      end
      test_b1_S366: begin
        IMAGE_addr <= 350;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 25;
        test_state <= test_b1_S367;
      end
      test_b1_S367: begin
        IMAGE_addr <= 351;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S368;
      end
      test_b1_S368: begin
        IMAGE_addr <= 352;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S369;
      end
      test_b1_S369: begin
        IMAGE_addr <= 353;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S370;
      end
      test_b1_S370: begin
        IMAGE_addr <= 354;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S371;
      end
      test_b1_S371: begin
        IMAGE_addr <= 355;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S372;
      end
      test_b1_S372: begin
        IMAGE_addr <= 356;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 29;
        test_state <= test_b1_S373;
      end
      test_b1_S373: begin
        IMAGE_addr <= 357;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S374;
      end
      test_b1_S374: begin
        IMAGE_addr <= 358;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S375;
      end
      test_b1_S375: begin
        IMAGE_addr <= 359;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S376;
      end
      test_b1_S376: begin
        IMAGE_addr <= 360;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S377;
      end
      test_b1_S377: begin
        IMAGE_addr <= 361;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 25;
        test_state <= test_b1_S378;
      end
      test_b1_S378: begin
        IMAGE_addr <= 362;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S379;
      end
      test_b1_S379: begin
        IMAGE_addr <= 363;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S380;
      end
      test_b1_S380: begin
        IMAGE_addr <= 364;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S381;
      end
      test_b1_S381: begin
        IMAGE_addr <= 365;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S382;
      end
      test_b1_S382: begin
        IMAGE_addr <= 366;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 29;
        test_state <= test_b1_S383;
      end
      test_b1_S383: begin
        IMAGE_addr <= 367;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 122;
        test_state <= test_b1_S384;
      end
      test_b1_S384: begin
        IMAGE_addr <= 368;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 345;
        test_state <= test_b1_S385;
      end
      test_b1_S385: begin
        IMAGE_addr <= 369;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S386;
      end
      test_b1_S386: begin
        IMAGE_addr <= 370;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S387;
      end
      test_b1_S387: begin
        IMAGE_addr <= 371;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S388;
      end
      test_b1_S388: begin
        IMAGE_addr <= 372;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S389;
      end
      test_b1_S389: begin
        IMAGE_addr <= 373;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S390;
      end
      test_b1_S390: begin
        IMAGE_addr <= 374;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 10;
        test_state <= test_b1_S391;
      end
      test_b1_S391: begin
        IMAGE_addr <= 375;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 359;
        test_state <= test_b1_S392;
      end
      test_b1_S392: begin
        IMAGE_addr <= 376;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S393;
      end
      test_b1_S393: begin
        IMAGE_addr <= 377;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S394;
      end
      test_b1_S394: begin
        IMAGE_addr <= 378;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 189;
        test_state <= test_b1_S395;
      end
      test_b1_S395: begin
        IMAGE_addr <= 379;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 25;
        test_state <= test_b1_S396;
      end
      test_b1_S396: begin
        IMAGE_addr <= 380;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 359;
        test_state <= test_b1_S397;
      end
      test_b1_S397: begin
        IMAGE_addr <= 381;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8;
        test_state <= test_b1_S398;
      end
      test_b1_S398: begin
        IMAGE_addr <= 382;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 378;
        test_state <= test_b1_S399;
      end
      test_b1_S399: begin
        IMAGE_addr <= 383;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S400;
      end
      test_b1_S400: begin
        IMAGE_addr <= 384;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S401;
      end
      test_b1_S401: begin
        IMAGE_addr <= 385;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8;
        test_state <= test_b1_S402;
      end
      test_b1_S402: begin
        IMAGE_addr <= 386;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6324;
        test_state <= test_b1_S403;
      end
      test_b1_S403: begin
        IMAGE_addr <= 387;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 378;
        test_state <= test_b1_S404;
      end
      test_b1_S404: begin
        IMAGE_addr <= 388;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S405;
      end
      test_b1_S405: begin
        IMAGE_addr <= 389;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S406;
      end
      test_b1_S406: begin
        IMAGE_addr <= 390;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S407;
      end
      test_b1_S407: begin
        IMAGE_addr <= 391;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S408;
      end
      test_b1_S408: begin
        IMAGE_addr <= 392;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S409;
      end
      test_b1_S409: begin
        IMAGE_addr <= 393;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 385;
        test_state <= test_b1_S410;
      end
      test_b1_S410: begin
        IMAGE_addr <= 394;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S411;
      end
      test_b1_S411: begin
        IMAGE_addr <= 395;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S412;
      end
      test_b1_S412: begin
        IMAGE_addr <= 396;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 32;
        test_state <= test_b1_S413;
      end
      test_b1_S413: begin
        IMAGE_addr <= 397;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4294967295;
        test_state <= test_b1_S414;
      end
      test_b1_S414: begin
        IMAGE_addr <= 398;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4294967295;
        test_state <= test_b1_S415;
      end
      test_b1_S415: begin
        IMAGE_addr <= 399;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4294967295;
        test_state <= test_b1_S416;
      end
      test_b1_S416: begin
        IMAGE_addr <= 400;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S417;
      end
      test_b1_S417: begin
        IMAGE_addr <= 401;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S418;
      end
      test_b1_S418: begin
        IMAGE_addr <= 402;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S419;
      end
      test_b1_S419: begin
        IMAGE_addr <= 403;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6;
        test_state <= test_b1_S420;
      end
      test_b1_S420: begin
        IMAGE_addr <= 404;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S421;
      end
      test_b1_S421: begin
        IMAGE_addr <= 405;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S422;
      end
      test_b1_S422: begin
        IMAGE_addr <= 406;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S423;
      end
      test_b1_S423: begin
        IMAGE_addr <= 407;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S424;
      end
      test_b1_S424: begin
        IMAGE_addr <= 408;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S425;
      end
      test_b1_S425: begin
        IMAGE_addr <= 409;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S426;
      end
      test_b1_S426: begin
        IMAGE_addr <= 410;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S427;
      end
      test_b1_S427: begin
        IMAGE_addr <= 411;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S428;
      end
      test_b1_S428: begin
        IMAGE_addr <= 412;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S429;
      end
      test_b1_S429: begin
        IMAGE_addr <= 413;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 127;
        test_state <= test_b1_S430;
      end
      test_b1_S430: begin
        IMAGE_addr <= 414;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 12;
        test_state <= test_b1_S431;
      end
      test_b1_S431: begin
        IMAGE_addr <= 415;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 419;
        test_state <= test_b1_S432;
      end
      test_b1_S432: begin
        IMAGE_addr <= 416;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S433;
      end
      test_b1_S433: begin
        IMAGE_addr <= 417;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S434;
      end
      test_b1_S434: begin
        IMAGE_addr <= 418;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8;
        test_state <= test_b1_S435;
      end
      test_b1_S435: begin
        IMAGE_addr <= 419;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S436;
      end
      test_b1_S436: begin
        IMAGE_addr <= 420;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S437;
      end
      test_b1_S437: begin
        IMAGE_addr <= 421;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 13;
        test_state <= test_b1_S438;
      end
      test_b1_S438: begin
        IMAGE_addr <= 422;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 12;
        test_state <= test_b1_S439;
      end
      test_b1_S439: begin
        IMAGE_addr <= 423;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 427;
        test_state <= test_b1_S440;
      end
      test_b1_S440: begin
        IMAGE_addr <= 424;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S441;
      end
      test_b1_S441: begin
        IMAGE_addr <= 425;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S442;
      end
      test_b1_S442: begin
        IMAGE_addr <= 426;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 10;
        test_state <= test_b1_S443;
      end
      test_b1_S443: begin
        IMAGE_addr <= 427;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S444;
      end
      test_b1_S444: begin
        IMAGE_addr <= 428;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 397;
        test_state <= test_b1_S445;
      end
      test_b1_S445: begin
        IMAGE_addr <= 429;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S446;
      end
      test_b1_S446: begin
        IMAGE_addr <= 430;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 25;
        test_state <= test_b1_S447;
      end
      test_b1_S447: begin
        IMAGE_addr <= 431;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S448;
      end
      test_b1_S448: begin
        IMAGE_addr <= 432;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S449;
      end
      test_b1_S449: begin
        IMAGE_addr <= 433;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S450;
      end
      test_b1_S450: begin
        IMAGE_addr <= 434;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 10;
        test_state <= test_b1_S451;
      end
      test_b1_S451: begin
        IMAGE_addr <= 435;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 12;
        test_state <= test_b1_S452;
      end
      test_b1_S452: begin
        IMAGE_addr <= 436;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 440;
        test_state <= test_b1_S453;
      end
      test_b1_S453: begin
        IMAGE_addr <= 437;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S454;
      end
      test_b1_S454: begin
        IMAGE_addr <= 438;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S455;
      end
      test_b1_S455: begin
        IMAGE_addr <= 439;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 32;
        test_state <= test_b1_S456;
      end
      test_b1_S456: begin
        IMAGE_addr <= 440;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S457;
      end
      test_b1_S457: begin
        IMAGE_addr <= 441;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 399;
        test_state <= test_b1_S458;
      end
      test_b1_S458: begin
        IMAGE_addr <= 442;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S459;
      end
      test_b1_S459: begin
        IMAGE_addr <= 443;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 25;
        test_state <= test_b1_S460;
      end
      test_b1_S460: begin
        IMAGE_addr <= 444;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 52;
        test_state <= test_b1_S461;
      end
      test_b1_S461: begin
        IMAGE_addr <= 445;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S462;
      end
      test_b1_S462: begin
        IMAGE_addr <= 446;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S463;
      end
      test_b1_S463: begin
        IMAGE_addr <= 447;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S464;
      end
      test_b1_S464: begin
        IMAGE_addr <= 448;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 12;
        test_state <= test_b1_S465;
      end
      test_b1_S465: begin
        IMAGE_addr <= 449;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 453;
        test_state <= test_b1_S466;
      end
      test_b1_S466: begin
        IMAGE_addr <= 450;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S467;
      end
      test_b1_S467: begin
        IMAGE_addr <= 451;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S468;
      end
      test_b1_S468: begin
        IMAGE_addr <= 452;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 32;
        test_state <= test_b1_S469;
      end
      test_b1_S469: begin
        IMAGE_addr <= 453;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S470;
      end
      test_b1_S470: begin
        IMAGE_addr <= 454;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S471;
      end
      test_b1_S471: begin
        IMAGE_addr <= 455;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S472;
      end
      test_b1_S472: begin
        IMAGE_addr <= 456;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S473;
      end
      test_b1_S473: begin
        IMAGE_addr <= 457;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S474;
      end
      test_b1_S474: begin
        IMAGE_addr <= 458;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S475;
      end
      test_b1_S475: begin
        IMAGE_addr <= 459;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 29;
        test_state <= test_b1_S476;
      end
      test_b1_S476: begin
        IMAGE_addr <= 460;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 122;
        test_state <= test_b1_S477;
      end
      test_b1_S477: begin
        IMAGE_addr <= 461;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S478;
      end
      test_b1_S478: begin
        IMAGE_addr <= 462;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S479;
      end
      test_b1_S479: begin
        IMAGE_addr <= 463;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 28;
        test_state <= test_b1_S480;
      end
      test_b1_S480: begin
        IMAGE_addr <= 464;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S481;
      end
      test_b1_S481: begin
        IMAGE_addr <= 465;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S482;
      end
      test_b1_S482: begin
        IMAGE_addr <= 466;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S483;
      end
      test_b1_S483: begin
        IMAGE_addr <= 467;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S484;
      end
      test_b1_S484: begin
        IMAGE_addr <= 468;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 455;
        test_state <= test_b1_S485;
      end
      test_b1_S485: begin
        IMAGE_addr <= 469;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 407;
        test_state <= test_b1_S486;
      end
      test_b1_S486: begin
        IMAGE_addr <= 470;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 32;
        test_state <= test_b1_S487;
      end
      test_b1_S487: begin
        IMAGE_addr <= 471;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S488;
      end
      test_b1_S488: begin
        IMAGE_addr <= 472;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S489;
      end
      test_b1_S489: begin
        IMAGE_addr <= 473;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 13;
        test_state <= test_b1_S490;
      end
      test_b1_S490: begin
        IMAGE_addr <= 474;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 478;
        test_state <= test_b1_S491;
      end
      test_b1_S491: begin
        IMAGE_addr <= 475;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 411;
        test_state <= test_b1_S492;
      end
      test_b1_S492: begin
        IMAGE_addr <= 476;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S493;
      end
      test_b1_S493: begin
        IMAGE_addr <= 477;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S494;
      end
      test_b1_S494: begin
        IMAGE_addr <= 478;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S495;
      end
      test_b1_S495: begin
        IMAGE_addr <= 479;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8;
        test_state <= test_b1_S496;
      end
      test_b1_S496: begin
        IMAGE_addr <= 480;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 468;
        test_state <= test_b1_S497;
      end
      test_b1_S497: begin
        IMAGE_addr <= 481;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S498;
      end
      test_b1_S498: begin
        IMAGE_addr <= 482;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S499;
      end
      test_b1_S499: begin
        IMAGE_addr <= 483;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S500;
      end
      test_b1_S500: begin
        IMAGE_addr <= 484;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S501;
      end
      test_b1_S501: begin
        IMAGE_addr <= 485;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8;
        test_state <= test_b1_S502;
      end
      test_b1_S502: begin
        IMAGE_addr <= 486;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 12;
        test_state <= test_b1_S503;
      end
      test_b1_S503: begin
        IMAGE_addr <= 487;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 494;
        test_state <= test_b1_S504;
      end
      test_b1_S504: begin
        IMAGE_addr <= 488;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S505;
      end
      test_b1_S505: begin
        IMAGE_addr <= 489;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S506;
      end
      test_b1_S506: begin
        IMAGE_addr <= 490;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 396;
        test_state <= test_b1_S507;
      end
      test_b1_S507: begin
        IMAGE_addr <= 491;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S508;
      end
      test_b1_S508: begin
        IMAGE_addr <= 492;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S509;
      end
      test_b1_S509: begin
        IMAGE_addr <= 493;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S510;
      end
      test_b1_S510: begin
        IMAGE_addr <= 494;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S511;
      end
      test_b1_S511: begin
        IMAGE_addr <= 495;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 359;
        test_state <= test_b1_S512;
      end
      test_b1_S512: begin
        IMAGE_addr <= 496;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S513;
      end
      test_b1_S513: begin
        IMAGE_addr <= 497;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S514;
      end
      test_b1_S514: begin
        IMAGE_addr <= 498;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S515;
      end
      test_b1_S515: begin
        IMAGE_addr <= 499;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 398;
        test_state <= test_b1_S516;
      end
      test_b1_S516: begin
        IMAGE_addr <= 500;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S517;
      end
      test_b1_S517: begin
        IMAGE_addr <= 501;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 25;
        test_state <= test_b1_S518;
      end
      test_b1_S518: begin
        IMAGE_addr <= 502;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 52;
        test_state <= test_b1_S519;
      end
      test_b1_S519: begin
        IMAGE_addr <= 503;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 466;
        test_state <= test_b1_S520;
      end
      test_b1_S520: begin
        IMAGE_addr <= 504;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 483;
        test_state <= test_b1_S521;
      end
      test_b1_S521: begin
        IMAGE_addr <= 505;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S522;
      end
      test_b1_S522: begin
        IMAGE_addr <= 506;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S523;
      end
      test_b1_S523: begin
        IMAGE_addr <= 507;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 396;
        test_state <= test_b1_S524;
      end
      test_b1_S524: begin
        IMAGE_addr <= 508;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S525;
      end
      test_b1_S525: begin
        IMAGE_addr <= 509;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 13;
        test_state <= test_b1_S526;
      end
      test_b1_S526: begin
        IMAGE_addr <= 510;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 515;
        test_state <= test_b1_S527;
      end
      test_b1_S527: begin
        IMAGE_addr <= 511;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S528;
      end
      test_b1_S528: begin
        IMAGE_addr <= 512;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 197;
        test_state <= test_b1_S529;
      end
      test_b1_S529: begin
        IMAGE_addr <= 513;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S530;
      end
      test_b1_S530: begin
        IMAGE_addr <= 514;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S531;
      end
      test_b1_S531: begin
        IMAGE_addr <= 515;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S532;
      end
      test_b1_S532: begin
        IMAGE_addr <= 516;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8;
        test_state <= test_b1_S533;
      end
      test_b1_S533: begin
        IMAGE_addr <= 517;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 503;
        test_state <= test_b1_S534;
      end
      test_b1_S534: begin
        IMAGE_addr <= 518;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S535;
      end
      test_b1_S535: begin
        IMAGE_addr <= 519;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S536;
      end
      test_b1_S536: begin
        IMAGE_addr <= 520;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S537;
      end
      test_b1_S537: begin
        IMAGE_addr <= 521;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 26;
        test_state <= test_b1_S538;
      end
      test_b1_S538: begin
        IMAGE_addr <= 522;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 400;
        test_state <= test_b1_S539;
      end
      test_b1_S539: begin
        IMAGE_addr <= 523;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 10;
        test_state <= test_b1_S540;
      end
      test_b1_S540: begin
        IMAGE_addr <= 524;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 529;
        test_state <= test_b1_S541;
      end
      test_b1_S541: begin
        IMAGE_addr <= 525;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S542;
      end
      test_b1_S542: begin
        IMAGE_addr <= 526;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 400;
        test_state <= test_b1_S543;
      end
      test_b1_S543: begin
        IMAGE_addr <= 527;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S544;
      end
      test_b1_S544: begin
        IMAGE_addr <= 528;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S545;
      end
      test_b1_S545: begin
        IMAGE_addr <= 529;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S546;
      end
      test_b1_S546: begin
        IMAGE_addr <= 530;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8;
        test_state <= test_b1_S547;
      end
      test_b1_S547: begin
        IMAGE_addr <= 531;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 359;
        test_state <= test_b1_S548;
      end
      test_b1_S548: begin
        IMAGE_addr <= 532;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S549;
      end
      test_b1_S549: begin
        IMAGE_addr <= 533;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S550;
      end
      test_b1_S550: begin
        IMAGE_addr <= 534;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 466;
        test_state <= test_b1_S551;
      end
      test_b1_S551: begin
        IMAGE_addr <= 535;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S552;
      end
      test_b1_S552: begin
        IMAGE_addr <= 536;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S553;
      end
      test_b1_S553: begin
        IMAGE_addr <= 537;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8;
        test_state <= test_b1_S554;
      end
      test_b1_S554: begin
        IMAGE_addr <= 538;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 12;
        test_state <= test_b1_S555;
      end
      test_b1_S555: begin
        IMAGE_addr <= 539;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 545;
        test_state <= test_b1_S556;
      end
      test_b1_S556: begin
        IMAGE_addr <= 540;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S557;
      end
      test_b1_S557: begin
        IMAGE_addr <= 541;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 27;
        test_state <= test_b1_S558;
      end
      test_b1_S558: begin
        IMAGE_addr <= 542;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 520;
        test_state <= test_b1_S559;
      end
      test_b1_S559: begin
        IMAGE_addr <= 543;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8;
        test_state <= test_b1_S560;
      end
      test_b1_S560: begin
        IMAGE_addr <= 544;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 534;
        test_state <= test_b1_S561;
      end
      test_b1_S561: begin
        IMAGE_addr <= 545;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S562;
      end
      test_b1_S562: begin
        IMAGE_addr <= 546;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 359;
        test_state <= test_b1_S563;
      end
      test_b1_S563: begin
        IMAGE_addr <= 547;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S564;
      end
      test_b1_S564: begin
        IMAGE_addr <= 548;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S565;
      end
      test_b1_S565: begin
        IMAGE_addr <= 549;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 396;
        test_state <= test_b1_S566;
      end
      test_b1_S566: begin
        IMAGE_addr <= 550;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S567;
      end
      test_b1_S567: begin
        IMAGE_addr <= 551;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 12;
        test_state <= test_b1_S568;
      end
      test_b1_S568: begin
        IMAGE_addr <= 552;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 556;
        test_state <= test_b1_S569;
      end
      test_b1_S569: begin
        IMAGE_addr <= 553;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S570;
      end
      test_b1_S570: begin
        IMAGE_addr <= 554;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S571;
      end
      test_b1_S571: begin
        IMAGE_addr <= 555;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S572;
      end
      test_b1_S572: begin
        IMAGE_addr <= 556;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S573;
      end
      test_b1_S573: begin
        IMAGE_addr <= 557;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 197;
        test_state <= test_b1_S574;
      end
      test_b1_S574: begin
        IMAGE_addr <= 558;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8;
        test_state <= test_b1_S575;
      end
      test_b1_S575: begin
        IMAGE_addr <= 559;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 534;
        test_state <= test_b1_S576;
      end
      test_b1_S576: begin
        IMAGE_addr <= 560;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S577;
      end
      test_b1_S577: begin
        IMAGE_addr <= 561;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S578;
      end
      test_b1_S578: begin
        IMAGE_addr <= 562;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S579;
      end
      test_b1_S579: begin
        IMAGE_addr <= 563;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S580;
      end
      test_b1_S580: begin
        IMAGE_addr <= 564;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S581;
      end
      test_b1_S581: begin
        IMAGE_addr <= 565;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 396;
        test_state <= test_b1_S582;
      end
      test_b1_S582: begin
        IMAGE_addr <= 566;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S583;
      end
      test_b1_S583: begin
        IMAGE_addr <= 567;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 400;
        test_state <= test_b1_S584;
      end
      test_b1_S584: begin
        IMAGE_addr <= 568;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 498;
        test_state <= test_b1_S585;
      end
      test_b1_S585: begin
        IMAGE_addr <= 569;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 534;
        test_state <= test_b1_S586;
      end
      test_b1_S586: begin
        IMAGE_addr <= 570;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S587;
      end
      test_b1_S587: begin
        IMAGE_addr <= 571;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S588;
      end
      test_b1_S588: begin
        IMAGE_addr <= 572;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S589;
      end
      test_b1_S589: begin
        IMAGE_addr <= 573;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 197;
        test_state <= test_b1_S590;
      end
      test_b1_S590: begin
        IMAGE_addr <= 574;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S591;
      end
      test_b1_S591: begin
        IMAGE_addr <= 575;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S592;
      end
      test_b1_S592: begin
        IMAGE_addr <= 576;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S593;
      end
      test_b1_S593: begin
        IMAGE_addr <= 577;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4294967295;
        test_state <= test_b1_S594;
      end
      test_b1_S594: begin
        IMAGE_addr <= 578;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S595;
      end
      test_b1_S595: begin
        IMAGE_addr <= 579;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S596;
      end
      test_b1_S596: begin
        IMAGE_addr <= 580;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 26;
        test_state <= test_b1_S597;
      end
      test_b1_S597: begin
        IMAGE_addr <= 581;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S598;
      end
      test_b1_S598: begin
        IMAGE_addr <= 582;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S599;
      end
      test_b1_S599: begin
        IMAGE_addr <= 583;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S600;
      end
      test_b1_S600: begin
        IMAGE_addr <= 584;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S601;
      end
      test_b1_S601: begin
        IMAGE_addr <= 585;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 26;
        test_state <= test_b1_S602;
      end
      test_b1_S602: begin
        IMAGE_addr <= 586;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 26;
        test_state <= test_b1_S603;
      end
      test_b1_S603: begin
        IMAGE_addr <= 587;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S604;
      end
      test_b1_S604: begin
        IMAGE_addr <= 588;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S605;
      end
      test_b1_S605: begin
        IMAGE_addr <= 589;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S606;
      end
      test_b1_S606: begin
        IMAGE_addr <= 590;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S607;
      end
      test_b1_S607: begin
        IMAGE_addr <= 591;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 26;
        test_state <= test_b1_S608;
      end
      test_b1_S608: begin
        IMAGE_addr <= 592;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 26;
        test_state <= test_b1_S609;
      end
      test_b1_S609: begin
        IMAGE_addr <= 593;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 26;
        test_state <= test_b1_S610;
      end
      test_b1_S610: begin
        IMAGE_addr <= 594;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S611;
      end
      test_b1_S611: begin
        IMAGE_addr <= 595;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S612;
      end
      test_b1_S612: begin
        IMAGE_addr <= 596;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S613;
      end
      test_b1_S613: begin
        IMAGE_addr <= 597;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S614;
      end
      test_b1_S614: begin
        IMAGE_addr <= 598;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5;
        test_state <= test_b1_S615;
      end
      test_b1_S615: begin
        IMAGE_addr <= 599;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 206;
        test_state <= test_b1_S616;
      end
      test_b1_S616: begin
        IMAGE_addr <= 600;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S617;
      end
      test_b1_S617: begin
        IMAGE_addr <= 601;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S618;
      end
      test_b1_S618: begin
        IMAGE_addr <= 602;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S619;
      end
      test_b1_S619: begin
        IMAGE_addr <= 603;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 213;
        test_state <= test_b1_S620;
      end
      test_b1_S620: begin
        IMAGE_addr <= 604;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S621;
      end
      test_b1_S621: begin
        IMAGE_addr <= 605;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S622;
      end
      test_b1_S622: begin
        IMAGE_addr <= 606;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S623;
      end
      test_b1_S623: begin
        IMAGE_addr <= 607;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S624;
      end
      test_b1_S624: begin
        IMAGE_addr <= 608;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 310;
        test_state <= test_b1_S625;
      end
      test_b1_S625: begin
        IMAGE_addr <= 609;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 213;
        test_state <= test_b1_S626;
      end
      test_b1_S626: begin
        IMAGE_addr <= 610;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 206;
        test_state <= test_b1_S627;
      end
      test_b1_S627: begin
        IMAGE_addr <= 611;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S628;
      end
      test_b1_S628: begin
        IMAGE_addr <= 612;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S629;
      end
      test_b1_S629: begin
        IMAGE_addr <= 613;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 213;
        test_state <= test_b1_S630;
      end
      test_b1_S630: begin
        IMAGE_addr <= 614;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6;
        test_state <= test_b1_S631;
      end
      test_b1_S631: begin
        IMAGE_addr <= 615;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 245;
        test_state <= test_b1_S632;
      end
      test_b1_S632: begin
        IMAGE_addr <= 616;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 206;
        test_state <= test_b1_S633;
      end
      test_b1_S633: begin
        IMAGE_addr <= 617;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S634;
      end
      test_b1_S634: begin
        IMAGE_addr <= 618;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S635;
      end
      test_b1_S635: begin
        IMAGE_addr <= 619;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S636;
      end
      test_b1_S636: begin
        IMAGE_addr <= 620;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S637;
      end
      test_b1_S637: begin
        IMAGE_addr <= 621;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S638;
      end
      test_b1_S638: begin
        IMAGE_addr <= 622;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S639;
      end
      test_b1_S639: begin
        IMAGE_addr <= 623;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S640;
      end
      test_b1_S640: begin
        IMAGE_addr <= 624;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 32;
        test_state <= test_b1_S641;
      end
      test_b1_S641: begin
        IMAGE_addr <= 625;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 562;
        test_state <= test_b1_S642;
      end
      test_b1_S642: begin
        IMAGE_addr <= 626;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 400;
        test_state <= test_b1_S643;
      end
      test_b1_S643: begin
        IMAGE_addr <= 627;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 596;
        test_state <= test_b1_S644;
      end
      test_b1_S644: begin
        IMAGE_addr <= 628;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S645;
      end
      test_b1_S645: begin
        IMAGE_addr <= 629;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S646;
      end
      test_b1_S646: begin
        IMAGE_addr <= 630;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S647;
      end
      test_b1_S647: begin
        IMAGE_addr <= 631;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S648;
      end
      test_b1_S648: begin
        IMAGE_addr <= 632;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S649;
      end
      test_b1_S649: begin
        IMAGE_addr <= 633;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S650;
      end
      test_b1_S650: begin
        IMAGE_addr <= 634;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 155;
        test_state <= test_b1_S651;
      end
      test_b1_S651: begin
        IMAGE_addr <= 635;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S652;
      end
      test_b1_S652: begin
        IMAGE_addr <= 636;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S653;
      end
      test_b1_S653: begin
        IMAGE_addr <= 637;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S654;
      end
      test_b1_S654: begin
        IMAGE_addr <= 638;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S655;
      end
      test_b1_S655: begin
        IMAGE_addr <= 639;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S656;
      end
      test_b1_S656: begin
        IMAGE_addr <= 640;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S657;
      end
      test_b1_S657: begin
        IMAGE_addr <= 641;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 147;
        test_state <= test_b1_S658;
      end
      test_b1_S658: begin
        IMAGE_addr <= 642;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S659;
      end
      test_b1_S659: begin
        IMAGE_addr <= 643;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S660;
      end
      test_b1_S660: begin
        IMAGE_addr <= 644;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S661;
      end
      test_b1_S661: begin
        IMAGE_addr <= 645;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S662;
      end
      test_b1_S662: begin
        IMAGE_addr <= 646;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S663;
      end
      test_b1_S663: begin
        IMAGE_addr <= 647;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 577;
        test_state <= test_b1_S664;
      end
      test_b1_S664: begin
        IMAGE_addr <= 648;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S665;
      end
      test_b1_S665: begin
        IMAGE_addr <= 649;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 25;
        test_state <= test_b1_S666;
      end
      test_b1_S666: begin
        IMAGE_addr <= 650;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S667;
      end
      test_b1_S667: begin
        IMAGE_addr <= 651;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S668;
      end
      test_b1_S668: begin
        IMAGE_addr <= 652;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S669;
      end
      test_b1_S669: begin
        IMAGE_addr <= 653;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 213;
        test_state <= test_b1_S670;
      end
      test_b1_S670: begin
        IMAGE_addr <= 654;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S671;
      end
      test_b1_S671: begin
        IMAGE_addr <= 655;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S672;
      end
      test_b1_S672: begin
        IMAGE_addr <= 656;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 213;
        test_state <= test_b1_S673;
      end
      test_b1_S673: begin
        IMAGE_addr <= 657;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S674;
      end
      test_b1_S674: begin
        IMAGE_addr <= 658;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S675;
      end
      test_b1_S675: begin
        IMAGE_addr <= 659;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S676;
      end
      test_b1_S676: begin
        IMAGE_addr <= 660;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S677;
      end
      test_b1_S677: begin
        IMAGE_addr <= 661;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 621;
        test_state <= test_b1_S678;
      end
      test_b1_S678: begin
        IMAGE_addr <= 662;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S679;
      end
      test_b1_S679: begin
        IMAGE_addr <= 663;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S680;
      end
      test_b1_S680: begin
        IMAGE_addr <= 664;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S681;
      end
      test_b1_S681: begin
        IMAGE_addr <= 665;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S682;
      end
      test_b1_S682: begin
        IMAGE_addr <= 666;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S683;
      end
      test_b1_S683: begin
        IMAGE_addr <= 667;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 578;
        test_state <= test_b1_S684;
      end
      test_b1_S684: begin
        IMAGE_addr <= 668;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S685;
      end
      test_b1_S685: begin
        IMAGE_addr <= 669;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 637;
        test_state <= test_b1_S686;
      end
      test_b1_S686: begin
        IMAGE_addr <= 670;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 644;
        test_state <= test_b1_S687;
      end
      test_b1_S687: begin
        IMAGE_addr <= 671;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S688;
      end
      test_b1_S688: begin
        IMAGE_addr <= 672;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S689;
      end
      test_b1_S689: begin
        IMAGE_addr <= 673;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S690;
      end
      test_b1_S690: begin
        IMAGE_addr <= 674;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S691;
      end
      test_b1_S691: begin
        IMAGE_addr <= 675;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S692;
      end
      test_b1_S692: begin
        IMAGE_addr <= 676;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 41;
        test_state <= test_b1_S693;
      end
      test_b1_S693: begin
        IMAGE_addr <= 677;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 562;
        test_state <= test_b1_S694;
      end
      test_b1_S694: begin
        IMAGE_addr <= 678;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S695;
      end
      test_b1_S695: begin
        IMAGE_addr <= 679;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S696;
      end
      test_b1_S696: begin
        IMAGE_addr <= 680;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S697;
      end
      test_b1_S697: begin
        IMAGE_addr <= 681;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S698;
      end
      test_b1_S698: begin
        IMAGE_addr <= 682;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6;
        test_state <= test_b1_S699;
      end
      test_b1_S699: begin
        IMAGE_addr <= 683;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 26;
        test_state <= test_b1_S700;
      end
      test_b1_S700: begin
        IMAGE_addr <= 684;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S701;
      end
      test_b1_S701: begin
        IMAGE_addr <= 685;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S702;
      end
      test_b1_S702: begin
        IMAGE_addr <= 686;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 27;
        test_state <= test_b1_S703;
      end
      test_b1_S703: begin
        IMAGE_addr <= 687;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5;
        test_state <= test_b1_S704;
      end
      test_b1_S704: begin
        IMAGE_addr <= 688;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 26;
        test_state <= test_b1_S705;
      end
      test_b1_S705: begin
        IMAGE_addr <= 689;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S706;
      end
      test_b1_S706: begin
        IMAGE_addr <= 690;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S707;
      end
      test_b1_S707: begin
        IMAGE_addr <= 691;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S708;
      end
      test_b1_S708: begin
        IMAGE_addr <= 692;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S709;
      end
      test_b1_S709: begin
        IMAGE_addr <= 693;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S710;
      end
      test_b1_S710: begin
        IMAGE_addr <= 694;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S711;
      end
      test_b1_S711: begin
        IMAGE_addr <= 695;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 213;
        test_state <= test_b1_S712;
      end
      test_b1_S712: begin
        IMAGE_addr <= 696;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 206;
        test_state <= test_b1_S713;
      end
      test_b1_S713: begin
        IMAGE_addr <= 697;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S714;
      end
      test_b1_S714: begin
        IMAGE_addr <= 698;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S715;
      end
      test_b1_S715: begin
        IMAGE_addr <= 699;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 213;
        test_state <= test_b1_S716;
      end
      test_b1_S716: begin
        IMAGE_addr <= 700;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S717;
      end
      test_b1_S717: begin
        IMAGE_addr <= 701;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S718;
      end
      test_b1_S718: begin
        IMAGE_addr <= 702;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S719;
      end
      test_b1_S719: begin
        IMAGE_addr <= 703;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S720;
      end
      test_b1_S720: begin
        IMAGE_addr <= 704;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S721;
      end
      test_b1_S721: begin
        IMAGE_addr <= 705;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 147;
        test_state <= test_b1_S722;
      end
      test_b1_S722: begin
        IMAGE_addr <= 706;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S723;
      end
      test_b1_S723: begin
        IMAGE_addr <= 707;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S724;
      end
      test_b1_S724: begin
        IMAGE_addr <= 708;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S725;
      end
      test_b1_S725: begin
        IMAGE_addr <= 709;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S726;
      end
      test_b1_S726: begin
        IMAGE_addr <= 710;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 222;
        test_state <= test_b1_S727;
      end
      test_b1_S727: begin
        IMAGE_addr <= 711;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S728;
      end
      test_b1_S728: begin
        IMAGE_addr <= 712;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S729;
      end
      test_b1_S729: begin
        IMAGE_addr <= 713;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S730;
      end
      test_b1_S730: begin
        IMAGE_addr <= 714;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 206;
        test_state <= test_b1_S731;
      end
      test_b1_S731: begin
        IMAGE_addr <= 715;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 132;
        test_state <= test_b1_S732;
      end
      test_b1_S732: begin
        IMAGE_addr <= 716;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S733;
      end
      test_b1_S733: begin
        IMAGE_addr <= 717;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S734;
      end
      test_b1_S734: begin
        IMAGE_addr <= 718;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S735;
      end
      test_b1_S735: begin
        IMAGE_addr <= 719;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S736;
      end
      test_b1_S736: begin
        IMAGE_addr <= 720;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S737;
      end
      test_b1_S737: begin
        IMAGE_addr <= 721;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S738;
      end
      test_b1_S738: begin
        IMAGE_addr <= 722;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 12;
        test_state <= test_b1_S739;
      end
      test_b1_S739: begin
        IMAGE_addr <= 723;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 727;
        test_state <= test_b1_S740;
      end
      test_b1_S740: begin
        IMAGE_addr <= 724;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 26;
        test_state <= test_b1_S741;
      end
      test_b1_S741: begin
        IMAGE_addr <= 725;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S742;
      end
      test_b1_S742: begin
        IMAGE_addr <= 726;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S743;
      end
      test_b1_S743: begin
        IMAGE_addr <= 727;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S744;
      end
      test_b1_S744: begin
        IMAGE_addr <= 728;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S745;
      end
      test_b1_S745: begin
        IMAGE_addr <= 729;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S746;
      end
      test_b1_S746: begin
        IMAGE_addr <= 730;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S747;
      end
      test_b1_S747: begin
        IMAGE_addr <= 731;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S748;
      end
      test_b1_S748: begin
        IMAGE_addr <= 732;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S749;
      end
      test_b1_S749: begin
        IMAGE_addr <= 733;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S750;
      end
      test_b1_S750: begin
        IMAGE_addr <= 734;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5;
        test_state <= test_b1_S751;
      end
      test_b1_S751: begin
        IMAGE_addr <= 735;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S752;
      end
      test_b1_S752: begin
        IMAGE_addr <= 736;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6;
        test_state <= test_b1_S753;
      end
      test_b1_S753: begin
        IMAGE_addr <= 737;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S754;
      end
      test_b1_S754: begin
        IMAGE_addr <= 738;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S755;
      end
      test_b1_S755: begin
        IMAGE_addr <= 739;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S756;
      end
      test_b1_S756: begin
        IMAGE_addr <= 740;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 13;
        test_state <= test_b1_S757;
      end
      test_b1_S757: begin
        IMAGE_addr <= 741;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 746;
        test_state <= test_b1_S758;
      end
      test_b1_S758: begin
        IMAGE_addr <= 742;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S759;
      end
      test_b1_S759: begin
        IMAGE_addr <= 743;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 183;
        test_state <= test_b1_S760;
      end
      test_b1_S760: begin
        IMAGE_addr <= 744;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S761;
      end
      test_b1_S761: begin
        IMAGE_addr <= 745;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S762;
      end
      test_b1_S762: begin
        IMAGE_addr <= 746;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S763;
      end
      test_b1_S763: begin
        IMAGE_addr <= 747;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S764;
      end
      test_b1_S764: begin
        IMAGE_addr <= 748;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 183;
        test_state <= test_b1_S765;
      end
      test_b1_S765: begin
        IMAGE_addr <= 749;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S766;
      end
      test_b1_S766: begin
        IMAGE_addr <= 750;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S767;
      end
      test_b1_S767: begin
        IMAGE_addr <= 751;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S768;
      end
      test_b1_S768: begin
        IMAGE_addr <= 752;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S769;
      end
      test_b1_S769: begin
        IMAGE_addr <= 753;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S770;
      end
      test_b1_S770: begin
        IMAGE_addr <= 754;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 730;
        test_state <= test_b1_S771;
      end
      test_b1_S771: begin
        IMAGE_addr <= 755;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 732;
        test_state <= test_b1_S772;
      end
      test_b1_S772: begin
        IMAGE_addr <= 756;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S773;
      end
      test_b1_S773: begin
        IMAGE_addr <= 757;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S774;
      end
      test_b1_S774: begin
        IMAGE_addr <= 758;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S775;
      end
      test_b1_S775: begin
        IMAGE_addr <= 759;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S776;
      end
      test_b1_S776: begin
        IMAGE_addr <= 760;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S777;
      end
      test_b1_S777: begin
        IMAGE_addr <= 761;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 730;
        test_state <= test_b1_S778;
      end
      test_b1_S778: begin
        IMAGE_addr <= 762;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S779;
      end
      test_b1_S779: begin
        IMAGE_addr <= 763;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 732;
        test_state <= test_b1_S780;
      end
      test_b1_S780: begin
        IMAGE_addr <= 764;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S781;
      end
      test_b1_S781: begin
        IMAGE_addr <= 765;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S782;
      end
      test_b1_S782: begin
        IMAGE_addr <= 766;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S783;
      end
      test_b1_S783: begin
        IMAGE_addr <= 767;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S784;
      end
      test_b1_S784: begin
        IMAGE_addr <= 768;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S785;
      end
      test_b1_S785: begin
        IMAGE_addr <= 769;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5;
        test_state <= test_b1_S786;
      end
      test_b1_S786: begin
        IMAGE_addr <= 770;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 183;
        test_state <= test_b1_S787;
      end
      test_b1_S787: begin
        IMAGE_addr <= 771;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6;
        test_state <= test_b1_S788;
      end
      test_b1_S788: begin
        IMAGE_addr <= 772;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S789;
      end
      test_b1_S789: begin
        IMAGE_addr <= 773;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S790;
      end
      test_b1_S790: begin
        IMAGE_addr <= 774;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S791;
      end
      test_b1_S791: begin
        IMAGE_addr <= 775;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S792;
      end
      test_b1_S792: begin
        IMAGE_addr <= 776;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 132;
        test_state <= test_b1_S793;
      end
      test_b1_S793: begin
        IMAGE_addr <= 777;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S794;
      end
      test_b1_S794: begin
        IMAGE_addr <= 778;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 183;
        test_state <= test_b1_S795;
      end
      test_b1_S795: begin
        IMAGE_addr <= 779;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 766;
        test_state <= test_b1_S796;
      end
      test_b1_S796: begin
        IMAGE_addr <= 780;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S797;
      end
      test_b1_S797: begin
        IMAGE_addr <= 781;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S798;
      end
      test_b1_S798: begin
        IMAGE_addr <= 782;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S799;
      end
      test_b1_S799: begin
        IMAGE_addr <= 783;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S800;
      end
      test_b1_S800: begin
        IMAGE_addr <= 784;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S801;
      end
      test_b1_S801: begin
        IMAGE_addr <= 785;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S802;
      end
      test_b1_S802: begin
        IMAGE_addr <= 786;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S803;
      end
      test_b1_S803: begin
        IMAGE_addr <= 787;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4294967295;
        test_state <= test_b1_S804;
      end
      test_b1_S804: begin
        IMAGE_addr <= 788;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S805;
      end
      test_b1_S805: begin
        IMAGE_addr <= 789;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S806;
      end
      test_b1_S806: begin
        IMAGE_addr <= 790;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S807;
      end
      test_b1_S807: begin
        IMAGE_addr <= 791;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S808;
      end
      test_b1_S808: begin
        IMAGE_addr <= 792;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 12;
        test_state <= test_b1_S809;
      end
      test_b1_S809: begin
        IMAGE_addr <= 793;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 796;
        test_state <= test_b1_S810;
      end
      test_b1_S810: begin
        IMAGE_addr <= 794;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8;
        test_state <= test_b1_S811;
      end
      test_b1_S811: begin
        IMAGE_addr <= 795;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 786;
        test_state <= test_b1_S812;
      end
      test_b1_S812: begin
        IMAGE_addr <= 796;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8;
        test_state <= test_b1_S813;
      end
      test_b1_S813: begin
        IMAGE_addr <= 797;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 782;
        test_state <= test_b1_S814;
      end
      test_b1_S814: begin
        IMAGE_addr <= 798;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S815;
      end
      test_b1_S815: begin
        IMAGE_addr <= 799;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S816;
      end
      test_b1_S816: begin
        IMAGE_addr <= 800;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 13;
        test_state <= test_b1_S817;
      end
      test_b1_S817: begin
        IMAGE_addr <= 801;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 804;
        test_state <= test_b1_S818;
      end
      test_b1_S818: begin
        IMAGE_addr <= 802;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8;
        test_state <= test_b1_S819;
      end
      test_b1_S819: begin
        IMAGE_addr <= 803;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 786;
        test_state <= test_b1_S820;
      end
      test_b1_S820: begin
        IMAGE_addr <= 804;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8;
        test_state <= test_b1_S821;
      end
      test_b1_S821: begin
        IMAGE_addr <= 805;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 782;
        test_state <= test_b1_S822;
      end
      test_b1_S822: begin
        IMAGE_addr <= 806;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S823;
      end
      test_b1_S823: begin
        IMAGE_addr <= 807;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S824;
      end
      test_b1_S824: begin
        IMAGE_addr <= 808;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 11;
        test_state <= test_b1_S825;
      end
      test_b1_S825: begin
        IMAGE_addr <= 809;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 812;
        test_state <= test_b1_S826;
      end
      test_b1_S826: begin
        IMAGE_addr <= 810;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8;
        test_state <= test_b1_S827;
      end
      test_b1_S827: begin
        IMAGE_addr <= 811;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 786;
        test_state <= test_b1_S828;
      end
      test_b1_S828: begin
        IMAGE_addr <= 812;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8;
        test_state <= test_b1_S829;
      end
      test_b1_S829: begin
        IMAGE_addr <= 813;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 782;
        test_state <= test_b1_S830;
      end
      test_b1_S830: begin
        IMAGE_addr <= 814;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S831;
      end
      test_b1_S831: begin
        IMAGE_addr <= 815;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S832;
      end
      test_b1_S832: begin
        IMAGE_addr <= 816;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 10;
        test_state <= test_b1_S833;
      end
      test_b1_S833: begin
        IMAGE_addr <= 817;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 820;
        test_state <= test_b1_S834;
      end
      test_b1_S834: begin
        IMAGE_addr <= 818;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8;
        test_state <= test_b1_S835;
      end
      test_b1_S835: begin
        IMAGE_addr <= 819;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 786;
        test_state <= test_b1_S836;
      end
      test_b1_S836: begin
        IMAGE_addr <= 820;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8;
        test_state <= test_b1_S837;
      end
      test_b1_S837: begin
        IMAGE_addr <= 821;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 782;
        test_state <= test_b1_S838;
      end
      test_b1_S838: begin
        IMAGE_addr <= 822;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S839;
      end
      test_b1_S839: begin
        IMAGE_addr <= 823;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S840;
      end
      test_b1_S840: begin
        IMAGE_addr <= 824;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 11;
        test_state <= test_b1_S841;
      end
      test_b1_S841: begin
        IMAGE_addr <= 825;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 828;
        test_state <= test_b1_S842;
      end
      test_b1_S842: begin
        IMAGE_addr <= 826;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8;
        test_state <= test_b1_S843;
      end
      test_b1_S843: begin
        IMAGE_addr <= 827;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 782;
        test_state <= test_b1_S844;
      end
      test_b1_S844: begin
        IMAGE_addr <= 828;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8;
        test_state <= test_b1_S845;
      end
      test_b1_S845: begin
        IMAGE_addr <= 829;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 786;
        test_state <= test_b1_S846;
      end
      test_b1_S846: begin
        IMAGE_addr <= 830;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S847;
      end
      test_b1_S847: begin
        IMAGE_addr <= 831;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S848;
      end
      test_b1_S848: begin
        IMAGE_addr <= 832;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 10;
        test_state <= test_b1_S849;
      end
      test_b1_S849: begin
        IMAGE_addr <= 833;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 836;
        test_state <= test_b1_S850;
      end
      test_b1_S850: begin
        IMAGE_addr <= 834;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8;
        test_state <= test_b1_S851;
      end
      test_b1_S851: begin
        IMAGE_addr <= 835;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 782;
        test_state <= test_b1_S852;
      end
      test_b1_S852: begin
        IMAGE_addr <= 836;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8;
        test_state <= test_b1_S853;
      end
      test_b1_S853: begin
        IMAGE_addr <= 837;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 786;
        test_state <= test_b1_S854;
      end
      test_b1_S854: begin
        IMAGE_addr <= 838;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S855;
      end
      test_b1_S855: begin
        IMAGE_addr <= 839;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S856;
      end
      test_b1_S856: begin
        IMAGE_addr <= 840;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S857;
      end
      test_b1_S857: begin
        IMAGE_addr <= 841;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S858;
      end
      test_b1_S858: begin
        IMAGE_addr <= 842;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5;
        test_state <= test_b1_S859;
      end
      test_b1_S859: begin
        IMAGE_addr <= 843;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 26;
        test_state <= test_b1_S860;
      end
      test_b1_S860: begin
        IMAGE_addr <= 844;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S861;
      end
      test_b1_S861: begin
        IMAGE_addr <= 845;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S862;
      end
      test_b1_S862: begin
        IMAGE_addr <= 846;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S863;
      end
      test_b1_S863: begin
        IMAGE_addr <= 847;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5;
        test_state <= test_b1_S864;
      end
      test_b1_S864: begin
        IMAGE_addr <= 848;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 26;
        test_state <= test_b1_S865;
      end
      test_b1_S865: begin
        IMAGE_addr <= 849;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6;
        test_state <= test_b1_S866;
      end
      test_b1_S866: begin
        IMAGE_addr <= 850;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S867;
      end
      test_b1_S867: begin
        IMAGE_addr <= 851;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6;
        test_state <= test_b1_S868;
      end
      test_b1_S868: begin
        IMAGE_addr <= 852;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 13;
        test_state <= test_b1_S869;
      end
      test_b1_S869: begin
        IMAGE_addr <= 853;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 860;
        test_state <= test_b1_S870;
      end
      test_b1_S870: begin
        IMAGE_addr <= 854;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S871;
      end
      test_b1_S871: begin
        IMAGE_addr <= 855;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S872;
      end
      test_b1_S872: begin
        IMAGE_addr <= 856;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S873;
      end
      test_b1_S873: begin
        IMAGE_addr <= 857;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 22;
        test_state <= test_b1_S874;
      end
      test_b1_S874: begin
        IMAGE_addr <= 858;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S875;
      end
      test_b1_S875: begin
        IMAGE_addr <= 859;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S876;
      end
      test_b1_S876: begin
        IMAGE_addr <= 860;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S877;
      end
      test_b1_S877: begin
        IMAGE_addr <= 861;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S878;
      end
      test_b1_S878: begin
        IMAGE_addr <= 862;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 12;
        test_state <= test_b1_S879;
      end
      test_b1_S879: begin
        IMAGE_addr <= 863;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 840;
        test_state <= test_b1_S880;
      end
      test_b1_S880: begin
        IMAGE_addr <= 864;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S881;
      end
      test_b1_S881: begin
        IMAGE_addr <= 865;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S882;
      end
      test_b1_S882: begin
        IMAGE_addr <= 866;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S883;
      end
      test_b1_S883: begin
        IMAGE_addr <= 867;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4294967295;
        test_state <= test_b1_S884;
      end
      test_b1_S884: begin
        IMAGE_addr <= 868;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S885;
      end
      test_b1_S885: begin
        IMAGE_addr <= 869;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S886;
      end
      test_b1_S886: begin
        IMAGE_addr <= 870;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 189;
        test_state <= test_b1_S887;
      end
      test_b1_S887: begin
        IMAGE_addr <= 871;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 25;
        test_state <= test_b1_S888;
      end
      test_b1_S888: begin
        IMAGE_addr <= 872;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S889;
      end
      test_b1_S889: begin
        IMAGE_addr <= 873;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8;
        test_state <= test_b1_S890;
      end
      test_b1_S890: begin
        IMAGE_addr <= 874;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 870;
        test_state <= test_b1_S891;
      end
      test_b1_S891: begin
        IMAGE_addr <= 875;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S892;
      end
      test_b1_S892: begin
        IMAGE_addr <= 876;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S893;
      end
      test_b1_S893: begin
        IMAGE_addr <= 877;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S894;
      end
      test_b1_S894: begin
        IMAGE_addr <= 878;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S895;
      end
      test_b1_S895: begin
        IMAGE_addr <= 879;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S896;
      end
      test_b1_S896: begin
        IMAGE_addr <= 880;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 870;
        test_state <= test_b1_S897;
      end
      test_b1_S897: begin
        IMAGE_addr <= 881;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 27;
        test_state <= test_b1_S898;
      end
      test_b1_S898: begin
        IMAGE_addr <= 882;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S899;
      end
      test_b1_S899: begin
        IMAGE_addr <= 883;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 17;
        test_state <= test_b1_S900;
      end
      test_b1_S900: begin
        IMAGE_addr <= 884;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S901;
      end
      test_b1_S901: begin
        IMAGE_addr <= 885;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S902;
      end
      test_b1_S902: begin
        IMAGE_addr <= 886;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S903;
      end
      test_b1_S903: begin
        IMAGE_addr <= 887;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S904;
      end
      test_b1_S904: begin
        IMAGE_addr <= 888;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S905;
      end
      test_b1_S905: begin
        IMAGE_addr <= 889;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 877;
        test_state <= test_b1_S906;
      end
      test_b1_S906: begin
        IMAGE_addr <= 890;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S907;
      end
      test_b1_S907: begin
        IMAGE_addr <= 891;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S908;
      end
      test_b1_S908: begin
        IMAGE_addr <= 892;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S909;
      end
      test_b1_S909: begin
        IMAGE_addr <= 893;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S910;
      end
      test_b1_S910: begin
        IMAGE_addr <= 894;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 886;
        test_state <= test_b1_S911;
      end
      test_b1_S911: begin
        IMAGE_addr <= 895;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S912;
      end
      test_b1_S912: begin
        IMAGE_addr <= 896;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S913;
      end
      test_b1_S913: begin
        IMAGE_addr <= 897;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 16;
        test_state <= test_b1_S914;
      end
      test_b1_S914: begin
        IMAGE_addr <= 898;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 206;
        test_state <= test_b1_S915;
      end
      test_b1_S915: begin
        IMAGE_addr <= 899;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 16;
        test_state <= test_b1_S916;
      end
      test_b1_S916: begin
        IMAGE_addr <= 900;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S917;
      end
      test_b1_S917: begin
        IMAGE_addr <= 901;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8;
        test_state <= test_b1_S918;
      end
      test_b1_S918: begin
        IMAGE_addr <= 902;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 213;
        test_state <= test_b1_S919;
      end
      test_b1_S919: begin
        IMAGE_addr <= 903;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 213;
        test_state <= test_b1_S920;
      end
      test_b1_S920: begin
        IMAGE_addr <= 904;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 206;
        test_state <= test_b1_S921;
      end
      test_b1_S921: begin
        IMAGE_addr <= 905;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S922;
      end
      test_b1_S922: begin
        IMAGE_addr <= 906;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 245;
        test_state <= test_b1_S923;
      end
      test_b1_S923: begin
        IMAGE_addr <= 907;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S924;
      end
      test_b1_S924: begin
        IMAGE_addr <= 908;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S925;
      end
      test_b1_S925: begin
        IMAGE_addr <= 909;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S926;
      end
      test_b1_S926: begin
        IMAGE_addr <= 910;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S927;
      end
      test_b1_S927: begin
        IMAGE_addr <= 911;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S928;
      end
      test_b1_S928: begin
        IMAGE_addr <= 912;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 256;
        test_state <= test_b1_S929;
      end
      test_b1_S929: begin
        IMAGE_addr <= 913;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S930;
      end
      test_b1_S930: begin
        IMAGE_addr <= 914;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S931;
      end
      test_b1_S931: begin
        IMAGE_addr <= 915;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S932;
      end
      test_b1_S932: begin
        IMAGE_addr <= 916;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S933;
      end
      test_b1_S933: begin
        IMAGE_addr <= 917;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S934;
      end
      test_b1_S934: begin
        IMAGE_addr <= 918;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 12;
        test_state <= test_b1_S935;
      end
      test_b1_S935: begin
        IMAGE_addr <= 919;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S936;
      end
      test_b1_S936: begin
        IMAGE_addr <= 920;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S937;
      end
      test_b1_S937: begin
        IMAGE_addr <= 921;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S938;
      end
      test_b1_S938: begin
        IMAGE_addr <= 922;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4294967295;
        test_state <= test_b1_S939;
      end
      test_b1_S939: begin
        IMAGE_addr <= 923;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S940;
      end
      test_b1_S940: begin
        IMAGE_addr <= 924;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4294967295;
        test_state <= test_b1_S941;
      end
      test_b1_S941: begin
        IMAGE_addr <= 925;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 10;
        test_state <= test_b1_S942;
      end
      test_b1_S942: begin
        IMAGE_addr <= 926;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 48;
        test_state <= test_b1_S943;
      end
      test_b1_S943: begin
        IMAGE_addr <= 927;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 49;
        test_state <= test_b1_S944;
      end
      test_b1_S944: begin
        IMAGE_addr <= 928;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 50;
        test_state <= test_b1_S945;
      end
      test_b1_S945: begin
        IMAGE_addr <= 929;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 51;
        test_state <= test_b1_S946;
      end
      test_b1_S946: begin
        IMAGE_addr <= 930;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 52;
        test_state <= test_b1_S947;
      end
      test_b1_S947: begin
        IMAGE_addr <= 931;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 53;
        test_state <= test_b1_S948;
      end
      test_b1_S948: begin
        IMAGE_addr <= 932;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 54;
        test_state <= test_b1_S949;
      end
      test_b1_S949: begin
        IMAGE_addr <= 933;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 55;
        test_state <= test_b1_S950;
      end
      test_b1_S950: begin
        IMAGE_addr <= 934;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 56;
        test_state <= test_b1_S951;
      end
      test_b1_S951: begin
        IMAGE_addr <= 935;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 57;
        test_state <= test_b1_S952;
      end
      test_b1_S952: begin
        IMAGE_addr <= 936;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 65;
        test_state <= test_b1_S953;
      end
      test_b1_S953: begin
        IMAGE_addr <= 937;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 66;
        test_state <= test_b1_S954;
      end
      test_b1_S954: begin
        IMAGE_addr <= 938;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 67;
        test_state <= test_b1_S955;
      end
      test_b1_S955: begin
        IMAGE_addr <= 939;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 68;
        test_state <= test_b1_S956;
      end
      test_b1_S956: begin
        IMAGE_addr <= 940;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 69;
        test_state <= test_b1_S957;
      end
      test_b1_S957: begin
        IMAGE_addr <= 941;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 70;
        test_state <= test_b1_S958;
      end
      test_b1_S958: begin
        IMAGE_addr <= 942;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S959;
      end
      test_b1_S959: begin
        IMAGE_addr <= 943;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S960;
      end
      test_b1_S960: begin
        IMAGE_addr <= 944;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S961;
      end
      test_b1_S961: begin
        IMAGE_addr <= 945;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S962;
      end
      test_b1_S962: begin
        IMAGE_addr <= 946;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 926;
        test_state <= test_b1_S963;
      end
      test_b1_S963: begin
        IMAGE_addr <= 947;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S964;
      end
      test_b1_S964: begin
        IMAGE_addr <= 948;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S965;
      end
      test_b1_S965: begin
        IMAGE_addr <= 949;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 943;
        test_state <= test_b1_S966;
      end
      test_b1_S966: begin
        IMAGE_addr <= 950;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 16;
        test_state <= test_b1_S967;
      end
      test_b1_S967: begin
        IMAGE_addr <= 951;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S968;
      end
      test_b1_S968: begin
        IMAGE_addr <= 952;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 132;
        test_state <= test_b1_S969;
      end
      test_b1_S969: begin
        IMAGE_addr <= 953;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 12;
        test_state <= test_b1_S970;
      end
      test_b1_S970: begin
        IMAGE_addr <= 954;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 958;
        test_state <= test_b1_S971;
      end
      test_b1_S971: begin
        IMAGE_addr <= 955;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S972;
      end
      test_b1_S972: begin
        IMAGE_addr <= 956;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 922;
        test_state <= test_b1_S973;
      end
      test_b1_S973: begin
        IMAGE_addr <= 957;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 147;
        test_state <= test_b1_S974;
      end
      test_b1_S974: begin
        IMAGE_addr <= 958;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S975;
      end
      test_b1_S975: begin
        IMAGE_addr <= 959;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S976;
      end
      test_b1_S976: begin
        IMAGE_addr <= 960;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 42;
        test_state <= test_b1_S977;
      end
      test_b1_S977: begin
        IMAGE_addr <= 961;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S978;
      end
      test_b1_S978: begin
        IMAGE_addr <= 962;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5;
        test_state <= test_b1_S979;
      end
      test_b1_S979: begin
        IMAGE_addr <= 963;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 949;
        test_state <= test_b1_S980;
      end
      test_b1_S980: begin
        IMAGE_addr <= 964;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6;
        test_state <= test_b1_S981;
      end
      test_b1_S981: begin
        IMAGE_addr <= 965;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 25;
        test_state <= test_b1_S982;
      end
      test_b1_S982: begin
        IMAGE_addr <= 966;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 42;
        test_state <= test_b1_S983;
      end
      test_b1_S983: begin
        IMAGE_addr <= 967;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8;
        test_state <= test_b1_S984;
      end
      test_b1_S984: begin
        IMAGE_addr <= 968;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 961;
        test_state <= test_b1_S985;
      end
      test_b1_S985: begin
        IMAGE_addr <= 969;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S986;
      end
      test_b1_S986: begin
        IMAGE_addr <= 970;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S987;
      end
      test_b1_S987: begin
        IMAGE_addr <= 971;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S988;
      end
      test_b1_S988: begin
        IMAGE_addr <= 972;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 925;
        test_state <= test_b1_S989;
      end
      test_b1_S989: begin
        IMAGE_addr <= 973;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S990;
      end
      test_b1_S990: begin
        IMAGE_addr <= 974;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S991;
      end
      test_b1_S991: begin
        IMAGE_addr <= 975;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S992;
      end
      test_b1_S992: begin
        IMAGE_addr <= 976;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 16;
        test_state <= test_b1_S993;
      end
      test_b1_S993: begin
        IMAGE_addr <= 977;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 10;
        test_state <= test_b1_S994;
      end
      test_b1_S994: begin
        IMAGE_addr <= 978;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 982;
        test_state <= test_b1_S995;
      end
      test_b1_S995: begin
        IMAGE_addr <= 979;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 960;
        test_state <= test_b1_S996;
      end
      test_b1_S996: begin
        IMAGE_addr <= 980;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S997;
      end
      test_b1_S997: begin
        IMAGE_addr <= 981;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S998;
      end
      test_b1_S998: begin
        IMAGE_addr <= 982;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S999;
      end
      test_b1_S999: begin
        IMAGE_addr <= 983;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S1000;
      end
      test_b1_S1000: begin
        IMAGE_addr <= 984;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S1001;
      end
      test_b1_S1001: begin
        IMAGE_addr <= 985;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S1002;
      end
      test_b1_S1002: begin
        IMAGE_addr <= 986;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 922;
        test_state <= test_b1_S1003;
      end
      test_b1_S1003: begin
        IMAGE_addr <= 987;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 155;
        test_state <= test_b1_S1004;
      end
      test_b1_S1004: begin
        IMAGE_addr <= 988;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 971;
        test_state <= test_b1_S1005;
      end
      test_b1_S1005: begin
        IMAGE_addr <= 989;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S1006;
      end
      test_b1_S1006: begin
        IMAGE_addr <= 990;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S1007;
      end
      test_b1_S1007: begin
        IMAGE_addr <= 991;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 922;
        test_state <= test_b1_S1008;
      end
      test_b1_S1008: begin
        IMAGE_addr <= 992;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S1009;
      end
      test_b1_S1009: begin
        IMAGE_addr <= 993;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S1010;
      end
      test_b1_S1010: begin
        IMAGE_addr <= 994;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S1011;
      end
      test_b1_S1011: begin
        IMAGE_addr <= 995;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S1012;
      end
      test_b1_S1012: begin
        IMAGE_addr <= 996;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 48;
        test_state <= test_b1_S1013;
      end
      test_b1_S1013: begin
        IMAGE_addr <= 997;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 17;
        test_state <= test_b1_S1014;
      end
      test_b1_S1014: begin
        IMAGE_addr <= 998;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S1015;
      end
      test_b1_S1015: begin
        IMAGE_addr <= 999;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 925;
        test_state <= test_b1_S1016;
      end
      test_b1_S1016: begin
        IMAGE_addr <= 1000;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S1017;
      end
      test_b1_S1017: begin
        IMAGE_addr <= 1001;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S1018;
      end
      test_b1_S1018: begin
        IMAGE_addr <= 1002;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 16;
        test_state <= test_b1_S1019;
      end
      test_b1_S1019: begin
        IMAGE_addr <= 1003;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 12;
        test_state <= test_b1_S1020;
      end
      test_b1_S1020: begin
        IMAGE_addr <= 1004;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1013;
        test_state <= test_b1_S1021;
      end
      test_b1_S1021: begin
        IMAGE_addr <= 1005;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S1022;
      end
      test_b1_S1022: begin
        IMAGE_addr <= 1006;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S1023;
      end
      test_b1_S1023: begin
        IMAGE_addr <= 1007;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 16;
        test_state <= test_b1_S1024;
      end
      test_b1_S1024: begin
        IMAGE_addr <= 1008;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 11;
        test_state <= test_b1_S1025;
      end
      test_b1_S1025: begin
        IMAGE_addr <= 1009;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1013;
        test_state <= test_b1_S1026;
      end
      test_b1_S1026: begin
        IMAGE_addr <= 1010;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S1027;
      end
      test_b1_S1027: begin
        IMAGE_addr <= 1011;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7;
        test_state <= test_b1_S1028;
      end
      test_b1_S1028: begin
        IMAGE_addr <= 1012;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 17;
        test_state <= test_b1_S1029;
      end
      test_b1_S1029: begin
        IMAGE_addr <= 1013;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S1030;
      end
      test_b1_S1030: begin
        IMAGE_addr <= 1014;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S1031;
      end
      test_b1_S1031: begin
        IMAGE_addr <= 1015;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S1032;
      end
      test_b1_S1032: begin
        IMAGE_addr <= 1016;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S1033;
      end
      test_b1_S1033: begin
        IMAGE_addr <= 1017;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S1034;
      end
      test_b1_S1034: begin
        IMAGE_addr <= 1018;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 45;
        test_state <= test_b1_S1035;
      end
      test_b1_S1035: begin
        IMAGE_addr <= 1019;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 12;
        test_state <= test_b1_S1036;
      end
      test_b1_S1036: begin
        IMAGE_addr <= 1020;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1029;
        test_state <= test_b1_S1037;
      end
      test_b1_S1037: begin
        IMAGE_addr <= 1021;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S1038;
      end
      test_b1_S1038: begin
        IMAGE_addr <= 1022;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4294967295;
        test_state <= test_b1_S1039;
      end
      test_b1_S1039: begin
        IMAGE_addr <= 1023;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S1040;
      end
      test_b1_S1040: begin
        IMAGE_addr <= 1024;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 923;
        test_state <= test_b1_S1041;
      end
      test_b1_S1041: begin
        IMAGE_addr <= 1025;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S1042;
      end
      test_b1_S1042: begin
        IMAGE_addr <= 1026;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 26;
        test_state <= test_b1_S1043;
      end
      test_b1_S1043: begin
        IMAGE_addr <= 1027;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S1044;
      end
      test_b1_S1044: begin
        IMAGE_addr <= 1028;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S1045;
      end
      test_b1_S1045: begin
        IMAGE_addr <= 1029;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S1046;
      end
      test_b1_S1046: begin
        IMAGE_addr <= 1030;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S1047;
      end
      test_b1_S1047: begin
        IMAGE_addr <= 1031;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S1048;
      end
      test_b1_S1048: begin
        IMAGE_addr <= 1032;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 923;
        test_state <= test_b1_S1049;
      end
      test_b1_S1049: begin
        IMAGE_addr <= 1033;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S1050;
      end
      test_b1_S1050: begin
        IMAGE_addr <= 1034;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S1051;
      end
      test_b1_S1051: begin
        IMAGE_addr <= 1035;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S1052;
      end
      test_b1_S1052: begin
        IMAGE_addr <= 1036;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S1053;
      end
      test_b1_S1053: begin
        IMAGE_addr <= 1037;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S1054;
      end
      test_b1_S1054: begin
        IMAGE_addr <= 1038;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 25;
        test_state <= test_b1_S1055;
      end
      test_b1_S1055: begin
        IMAGE_addr <= 1039;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 995;
        test_state <= test_b1_S1056;
      end
      test_b1_S1056: begin
        IMAGE_addr <= 1040;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S1057;
      end
      test_b1_S1057: begin
        IMAGE_addr <= 1041;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 921;
        test_state <= test_b1_S1058;
      end
      test_b1_S1058: begin
        IMAGE_addr <= 1042;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S1059;
      end
      test_b1_S1059: begin
        IMAGE_addr <= 1043;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S1060;
      end
      test_b1_S1060: begin
        IMAGE_addr <= 1044;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 925;
        test_state <= test_b1_S1061;
      end
      test_b1_S1061: begin
        IMAGE_addr <= 1045;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S1062;
      end
      test_b1_S1062: begin
        IMAGE_addr <= 1046;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 18;
        test_state <= test_b1_S1063;
      end
      test_b1_S1063: begin
        IMAGE_addr <= 1047;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 16;
        test_state <= test_b1_S1064;
      end
      test_b1_S1064: begin
        IMAGE_addr <= 1048;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S1065;
      end
      test_b1_S1065: begin
        IMAGE_addr <= 1049;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 921;
        test_state <= test_b1_S1066;
      end
      test_b1_S1066: begin
        IMAGE_addr <= 1050;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S1067;
      end
      test_b1_S1067: begin
        IMAGE_addr <= 1051;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 26;
        test_state <= test_b1_S1068;
      end
      test_b1_S1068: begin
        IMAGE_addr <= 1052;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8;
        test_state <= test_b1_S1069;
      end
      test_b1_S1069: begin
        IMAGE_addr <= 1053;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1036;
        test_state <= test_b1_S1070;
      end
      test_b1_S1070: begin
        IMAGE_addr <= 1054;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S1071;
      end
      test_b1_S1071: begin
        IMAGE_addr <= 1055;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S1072;
      end
      test_b1_S1072: begin
        IMAGE_addr <= 1056;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1073;
      end
      test_b1_S1073: begin
        IMAGE_addr <= 1057;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1074;
      end
      test_b1_S1074: begin
        IMAGE_addr <= 1058;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1015;
        test_state <= test_b1_S1075;
      end
      test_b1_S1075: begin
        IMAGE_addr <= 1059;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S1076;
      end
      test_b1_S1076: begin
        IMAGE_addr <= 1060;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1077;
      end
      test_b1_S1077: begin
        IMAGE_addr <= 1061;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S1078;
      end
      test_b1_S1078: begin
        IMAGE_addr <= 1062;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 921;
        test_state <= test_b1_S1079;
      end
      test_b1_S1079: begin
        IMAGE_addr <= 1063;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S1080;
      end
      test_b1_S1080: begin
        IMAGE_addr <= 1064;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1036;
        test_state <= test_b1_S1081;
      end
      test_b1_S1081: begin
        IMAGE_addr <= 1065;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S1082;
      end
      test_b1_S1082: begin
        IMAGE_addr <= 1066;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S1083;
      end
      test_b1_S1083: begin
        IMAGE_addr <= 1067;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 921;
        test_state <= test_b1_S1084;
      end
      test_b1_S1084: begin
        IMAGE_addr <= 1068;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S1085;
      end
      test_b1_S1085: begin
        IMAGE_addr <= 1069;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S1086;
      end
      test_b1_S1086: begin
        IMAGE_addr <= 1070;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 923;
        test_state <= test_b1_S1087;
      end
      test_b1_S1087: begin
        IMAGE_addr <= 1071;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S1088;
      end
      test_b1_S1088: begin
        IMAGE_addr <= 1072;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 18;
        test_state <= test_b1_S1089;
      end
      test_b1_S1089: begin
        IMAGE_addr <= 1073;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S1090;
      end
      test_b1_S1090: begin
        IMAGE_addr <= 1074;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S1091;
      end
      test_b1_S1091: begin
        IMAGE_addr <= 1075;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S1092;
      end
      test_b1_S1092: begin
        IMAGE_addr <= 1076;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S1093;
      end
      test_b1_S1093: begin
        IMAGE_addr <= 1077;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 25;
        test_state <= test_b1_S1094;
      end
      test_b1_S1094: begin
        IMAGE_addr <= 1078;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 985;
        test_state <= test_b1_S1095;
      end
      test_b1_S1095: begin
        IMAGE_addr <= 1079;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S1096;
      end
      test_b1_S1096: begin
        IMAGE_addr <= 1080;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 924;
        test_state <= test_b1_S1097;
      end
      test_b1_S1097: begin
        IMAGE_addr <= 1081;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S1098;
      end
      test_b1_S1098: begin
        IMAGE_addr <= 1082;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 20;
        test_state <= test_b1_S1099;
      end
      test_b1_S1099: begin
        IMAGE_addr <= 1083;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S1100;
      end
      test_b1_S1100: begin
        IMAGE_addr <= 1084;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 924;
        test_state <= test_b1_S1101;
      end
      test_b1_S1101: begin
        IMAGE_addr <= 1085;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S1102;
      end
      test_b1_S1102: begin
        IMAGE_addr <= 1086;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 26;
        test_state <= test_b1_S1103;
      end
      test_b1_S1103: begin
        IMAGE_addr <= 1087;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8;
        test_state <= test_b1_S1104;
      end
      test_b1_S1104: begin
        IMAGE_addr <= 1088;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1075;
        test_state <= test_b1_S1105;
      end
      test_b1_S1105: begin
        IMAGE_addr <= 1089;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S1106;
      end
      test_b1_S1106: begin
        IMAGE_addr <= 1090;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S1107;
      end
      test_b1_S1107: begin
        IMAGE_addr <= 1091;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1108;
      end
      test_b1_S1108: begin
        IMAGE_addr <= 1092;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1109;
      end
      test_b1_S1109: begin
        IMAGE_addr <= 1093;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1015;
        test_state <= test_b1_S1110;
      end
      test_b1_S1110: begin
        IMAGE_addr <= 1094;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S1111;
      end
      test_b1_S1111: begin
        IMAGE_addr <= 1095;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 924;
        test_state <= test_b1_S1112;
      end
      test_b1_S1112: begin
        IMAGE_addr <= 1096;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 147;
        test_state <= test_b1_S1113;
      end
      test_b1_S1113: begin
        IMAGE_addr <= 1097;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1075;
        test_state <= test_b1_S1114;
      end
      test_b1_S1114: begin
        IMAGE_addr <= 1098;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S1115;
      end
      test_b1_S1115: begin
        IMAGE_addr <= 1099;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S1116;
      end
      test_b1_S1116: begin
        IMAGE_addr <= 1100;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 924;
        test_state <= test_b1_S1117;
      end
      test_b1_S1117: begin
        IMAGE_addr <= 1101;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S1118;
      end
      test_b1_S1118: begin
        IMAGE_addr <= 1102;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S1119;
      end
      test_b1_S1119: begin
        IMAGE_addr <= 1103;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S1120;
      end
      test_b1_S1120: begin
        IMAGE_addr <= 1104;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1000000;
        test_state <= test_b1_S1121;
      end
      test_b1_S1121: begin
        IMAGE_addr <= 1105;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1122;
      end
      test_b1_S1122: begin
        IMAGE_addr <= 1106;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1123;
      end
      test_b1_S1123: begin
        IMAGE_addr <= 1107;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1124;
      end
      test_b1_S1124: begin
        IMAGE_addr <= 1108;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 108;
        test_state <= test_b1_S1125;
      end
      test_b1_S1125: begin
        IMAGE_addr <= 1109;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 39;
        test_state <= test_b1_S1126;
      end
      test_b1_S1126: begin
        IMAGE_addr <= 1110;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1127;
      end
      test_b1_S1127: begin
        IMAGE_addr <= 1111;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1128;
      end
      test_b1_S1128: begin
        IMAGE_addr <= 1112;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S1129;
      end
      test_b1_S1129: begin
        IMAGE_addr <= 1113;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7;
        test_state <= test_b1_S1130;
      end
      test_b1_S1130: begin
        IMAGE_addr <= 1114;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 391;
        test_state <= test_b1_S1131;
      end
      test_b1_S1131: begin
        IMAGE_addr <= 1115;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S1132;
      end
      test_b1_S1132: begin
        IMAGE_addr <= 1116;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 32;
        test_state <= test_b1_S1133;
      end
      test_b1_S1133: begin
        IMAGE_addr <= 1117;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 359;
        test_state <= test_b1_S1134;
      end
      test_b1_S1134: begin
        IMAGE_addr <= 1118;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S1135;
      end
      test_b1_S1135: begin
        IMAGE_addr <= 1119;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 13;
        test_state <= test_b1_S1136;
      end
      test_b1_S1136: begin
        IMAGE_addr <= 1120;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 391;
        test_state <= test_b1_S1137;
      end
      test_b1_S1137: begin
        IMAGE_addr <= 1121;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S1138;
      end
      test_b1_S1138: begin
        IMAGE_addr <= 1122;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 32;
        test_state <= test_b1_S1139;
      end
      test_b1_S1139: begin
        IMAGE_addr <= 1123;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 359;
        test_state <= test_b1_S1140;
      end
      test_b1_S1140: begin
        IMAGE_addr <= 1124;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S1141;
      end
      test_b1_S1141: begin
        IMAGE_addr <= 1125;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 40;
        test_state <= test_b1_S1142;
      end
      test_b1_S1142: begin
        IMAGE_addr <= 1126;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 359;
        test_state <= test_b1_S1143;
      end
      test_b1_S1143: begin
        IMAGE_addr <= 1127;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S1144;
      end
      test_b1_S1144: begin
        IMAGE_addr <= 1128;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 18;
        test_state <= test_b1_S1145;
      end
      test_b1_S1145: begin
        IMAGE_addr <= 1129;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 391;
        test_state <= test_b1_S1146;
      end
      test_b1_S1146: begin
        IMAGE_addr <= 1130;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S1147;
      end
      test_b1_S1147: begin
        IMAGE_addr <= 1131;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 41;
        test_state <= test_b1_S1148;
      end
      test_b1_S1148: begin
        IMAGE_addr <= 1132;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 359;
        test_state <= test_b1_S1149;
      end
      test_b1_S1149: begin
        IMAGE_addr <= 1133;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 371;
        test_state <= test_b1_S1150;
      end
      test_b1_S1150: begin
        IMAGE_addr <= 1134;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S1151;
      end
      test_b1_S1151: begin
        IMAGE_addr <= 1135;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S1152;
      end
      test_b1_S1152: begin
        IMAGE_addr <= 1136;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S1153;
      end
      test_b1_S1153: begin
        IMAGE_addr <= 1137;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5;
        test_state <= test_b1_S1154;
      end
      test_b1_S1154: begin
        IMAGE_addr <= 1138;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 29;
        test_state <= test_b1_S1155;
      end
      test_b1_S1155: begin
        IMAGE_addr <= 1139;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 122;
        test_state <= test_b1_S1156;
      end
      test_b1_S1156: begin
        IMAGE_addr <= 1140;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S1157;
      end
      test_b1_S1157: begin
        IMAGE_addr <= 1141;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5;
        test_state <= test_b1_S1158;
      end
      test_b1_S1158: begin
        IMAGE_addr <= 1142;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 28;
        test_state <= test_b1_S1159;
      end
      test_b1_S1159: begin
        IMAGE_addr <= 1143;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S1160;
      end
      test_b1_S1160: begin
        IMAGE_addr <= 1144;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S1161;
      end
      test_b1_S1161: begin
        IMAGE_addr <= 1145;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S1162;
      end
      test_b1_S1162: begin
        IMAGE_addr <= 1146;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4294967295;
        test_state <= test_b1_S1163;
      end
      test_b1_S1163: begin
        IMAGE_addr <= 1147;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1136;
        test_state <= test_b1_S1164;
      end
      test_b1_S1164: begin
        IMAGE_addr <= 1148;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S1165;
      end
      test_b1_S1165: begin
        IMAGE_addr <= 1149;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1104;
        test_state <= test_b1_S1166;
      end
      test_b1_S1166: begin
        IMAGE_addr <= 1150;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S1167;
      end
      test_b1_S1167: begin
        IMAGE_addr <= 1151;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S1168;
      end
      test_b1_S1168: begin
        IMAGE_addr <= 1152;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4294967294;
        test_state <= test_b1_S1169;
      end
      test_b1_S1169: begin
        IMAGE_addr <= 1153;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1136;
        test_state <= test_b1_S1170;
      end
      test_b1_S1170: begin
        IMAGE_addr <= 1154;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S1171;
      end
      test_b1_S1171: begin
        IMAGE_addr <= 1155;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1105;
        test_state <= test_b1_S1172;
      end
      test_b1_S1172: begin
        IMAGE_addr <= 1156;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S1173;
      end
      test_b1_S1173: begin
        IMAGE_addr <= 1157;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S1174;
      end
      test_b1_S1174: begin
        IMAGE_addr <= 1158;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4294967293;
        test_state <= test_b1_S1175;
      end
      test_b1_S1175: begin
        IMAGE_addr <= 1159;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1136;
        test_state <= test_b1_S1176;
      end
      test_b1_S1176: begin
        IMAGE_addr <= 1160;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S1177;
      end
      test_b1_S1177: begin
        IMAGE_addr <= 1161;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1106;
        test_state <= test_b1_S1178;
      end
      test_b1_S1178: begin
        IMAGE_addr <= 1162;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S1179;
      end
      test_b1_S1179: begin
        IMAGE_addr <= 1163;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S1180;
      end
      test_b1_S1180: begin
        IMAGE_addr <= 1164;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4294967292;
        test_state <= test_b1_S1181;
      end
      test_b1_S1181: begin
        IMAGE_addr <= 1165;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1136;
        test_state <= test_b1_S1182;
      end
      test_b1_S1182: begin
        IMAGE_addr <= 1166;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S1183;
      end
      test_b1_S1183: begin
        IMAGE_addr <= 1167;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1107;
        test_state <= test_b1_S1184;
      end
      test_b1_S1184: begin
        IMAGE_addr <= 1168;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S1185;
      end
      test_b1_S1185: begin
        IMAGE_addr <= 1169;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S1186;
      end
      test_b1_S1186: begin
        IMAGE_addr <= 1170;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4294967285;
        test_state <= test_b1_S1187;
      end
      test_b1_S1187: begin
        IMAGE_addr <= 1171;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1136;
        test_state <= test_b1_S1188;
      end
      test_b1_S1188: begin
        IMAGE_addr <= 1172;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S1189;
      end
      test_b1_S1189: begin
        IMAGE_addr <= 1173;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1108;
        test_state <= test_b1_S1190;
      end
      test_b1_S1190: begin
        IMAGE_addr <= 1174;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S1191;
      end
      test_b1_S1191: begin
        IMAGE_addr <= 1175;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S1192;
      end
      test_b1_S1192: begin
        IMAGE_addr <= 1176;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4294967284;
        test_state <= test_b1_S1193;
      end
      test_b1_S1193: begin
        IMAGE_addr <= 1177;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1136;
        test_state <= test_b1_S1194;
      end
      test_b1_S1194: begin
        IMAGE_addr <= 1178;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S1195;
      end
      test_b1_S1195: begin
        IMAGE_addr <= 1179;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1109;
        test_state <= test_b1_S1196;
      end
      test_b1_S1196: begin
        IMAGE_addr <= 1180;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S1197;
      end
      test_b1_S1197: begin
        IMAGE_addr <= 1181;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1110;
        test_state <= test_b1_S1198;
      end
      test_b1_S1198: begin
        IMAGE_addr <= 1182;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S1199;
      end
      test_b1_S1199: begin
        IMAGE_addr <= 1183;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S1200;
      end
      test_b1_S1200: begin
        IMAGE_addr <= 1184;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2314;
        test_state <= test_b1_S1201;
      end
      test_b1_S1201: begin
        IMAGE_addr <= 1185;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4294967295;
        test_state <= test_b1_S1202;
      end
      test_b1_S1202: begin
        IMAGE_addr <= 1186;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S1203;
      end
      test_b1_S1203: begin
        IMAGE_addr <= 1187;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1185;
        test_state <= test_b1_S1204;
      end
      test_b1_S1204: begin
        IMAGE_addr <= 1188;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 155;
        test_state <= test_b1_S1205;
      end
      test_b1_S1205: begin
        IMAGE_addr <= 1189;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S1206;
      end
      test_b1_S1206: begin
        IMAGE_addr <= 1190;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1184;
        test_state <= test_b1_S1207;
      end
      test_b1_S1207: begin
        IMAGE_addr <= 1191;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S1208;
      end
      test_b1_S1208: begin
        IMAGE_addr <= 1192;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S1209;
      end
      test_b1_S1209: begin
        IMAGE_addr <= 1193;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S1210;
      end
      test_b1_S1210: begin
        IMAGE_addr <= 1194;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S1211;
      end
      test_b1_S1211: begin
        IMAGE_addr <= 1195;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S1212;
      end
      test_b1_S1212: begin
        IMAGE_addr <= 1196;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S1213;
      end
      test_b1_S1213: begin
        IMAGE_addr <= 1197;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S1214;
      end
      test_b1_S1214: begin
        IMAGE_addr <= 1198;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5;
        test_state <= test_b1_S1215;
      end
      test_b1_S1215: begin
        IMAGE_addr <= 1199;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S1216;
      end
      test_b1_S1216: begin
        IMAGE_addr <= 1200;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S1217;
      end
      test_b1_S1217: begin
        IMAGE_addr <= 1201;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1185;
        test_state <= test_b1_S1218;
      end
      test_b1_S1218: begin
        IMAGE_addr <= 1202;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S1219;
      end
      test_b1_S1219: begin
        IMAGE_addr <= 1203;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S1220;
      end
      test_b1_S1220: begin
        IMAGE_addr <= 1204;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S1221;
      end
      test_b1_S1221: begin
        IMAGE_addr <= 1205;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S1222;
      end
      test_b1_S1222: begin
        IMAGE_addr <= 1206;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 589;
        test_state <= test_b1_S1223;
      end
      test_b1_S1223: begin
        IMAGE_addr <= 1207;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S1224;
      end
      test_b1_S1224: begin
        IMAGE_addr <= 1208;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1184;
        test_state <= test_b1_S1225;
      end
      test_b1_S1225: begin
        IMAGE_addr <= 1209;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S1226;
      end
      test_b1_S1226: begin
        IMAGE_addr <= 1210;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 838;
        test_state <= test_b1_S1227;
      end
      test_b1_S1227: begin
        IMAGE_addr <= 1211;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S1228;
      end
      test_b1_S1228: begin
        IMAGE_addr <= 1212;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S1229;
      end
      test_b1_S1229: begin
        IMAGE_addr <= 1213;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1205;
        test_state <= test_b1_S1230;
      end
      test_b1_S1230: begin
        IMAGE_addr <= 1214;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S1231;
      end
      test_b1_S1231: begin
        IMAGE_addr <= 1215;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1232;
      end
      test_b1_S1232: begin
        IMAGE_addr <= 1216;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 13;
        test_state <= test_b1_S1233;
      end
      test_b1_S1233: begin
        IMAGE_addr <= 1217;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1226;
        test_state <= test_b1_S1234;
      end
      test_b1_S1234: begin
        IMAGE_addr <= 1218;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S1235;
      end
      test_b1_S1235: begin
        IMAGE_addr <= 1219;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5;
        test_state <= test_b1_S1236;
      end
      test_b1_S1236: begin
        IMAGE_addr <= 1220;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S1237;
      end
      test_b1_S1237: begin
        IMAGE_addr <= 1221;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S1238;
      end
      test_b1_S1238: begin
        IMAGE_addr <= 1222;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1185;
        test_state <= test_b1_S1239;
      end
      test_b1_S1239: begin
        IMAGE_addr <= 1223;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 147;
        test_state <= test_b1_S1240;
      end
      test_b1_S1240: begin
        IMAGE_addr <= 1224;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S1241;
      end
      test_b1_S1241: begin
        IMAGE_addr <= 1225;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S1242;
      end
      test_b1_S1242: begin
        IMAGE_addr <= 1226;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 72;
        test_state <= test_b1_S1243;
      end
      test_b1_S1243: begin
        IMAGE_addr <= 1227;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 25;
        test_state <= test_b1_S1244;
      end
      test_b1_S1244: begin
        IMAGE_addr <= 1228;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8;
        test_state <= test_b1_S1245;
      end
      test_b1_S1245: begin
        IMAGE_addr <= 1229;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1213;
        test_state <= test_b1_S1246;
      end
      test_b1_S1246: begin
        IMAGE_addr <= 1230;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S1247;
      end
      test_b1_S1247: begin
        IMAGE_addr <= 1231;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S1248;
      end
      test_b1_S1248: begin
        IMAGE_addr <= 1232;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8;
        test_state <= test_b1_S1249;
      end
      test_b1_S1249: begin
        IMAGE_addr <= 1233;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5452;
        test_state <= test_b1_S1250;
      end
      test_b1_S1250: begin
        IMAGE_addr <= 1234;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1186;
        test_state <= test_b1_S1251;
      end
      test_b1_S1251: begin
        IMAGE_addr <= 1235;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1213;
        test_state <= test_b1_S1252;
      end
      test_b1_S1252: begin
        IMAGE_addr <= 1236;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1197;
        test_state <= test_b1_S1253;
      end
      test_b1_S1253: begin
        IMAGE_addr <= 1237;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S1254;
      end
      test_b1_S1254: begin
        IMAGE_addr <= 1238;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S1255;
      end
      test_b1_S1255: begin
        IMAGE_addr <= 1239;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1256;
      end
      test_b1_S1256: begin
        IMAGE_addr <= 1240;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1257;
      end
      test_b1_S1257: begin
        IMAGE_addr <= 1241;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S1258;
      end
      test_b1_S1258: begin
        IMAGE_addr <= 1242;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 32;
        test_state <= test_b1_S1259;
      end
      test_b1_S1259: begin
        IMAGE_addr <= 1243;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 562;
        test_state <= test_b1_S1260;
      end
      test_b1_S1260: begin
        IMAGE_addr <= 1244;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 400;
        test_state <= test_b1_S1261;
      end
      test_b1_S1261: begin
        IMAGE_addr <= 1245;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1232;
        test_state <= test_b1_S1262;
      end
      test_b1_S1262: begin
        IMAGE_addr <= 1246;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S1263;
      end
      test_b1_S1263: begin
        IMAGE_addr <= 1247;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1264;
      end
      test_b1_S1264: begin
        IMAGE_addr <= 1248;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 13;
        test_state <= test_b1_S1265;
      end
      test_b1_S1265: begin
        IMAGE_addr <= 1249;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1254;
        test_state <= test_b1_S1266;
      end
      test_b1_S1266: begin
        IMAGE_addr <= 1250;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 583;
        test_state <= test_b1_S1267;
      end
      test_b1_S1267: begin
        IMAGE_addr <= 1251;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S1268;
      end
      test_b1_S1268: begin
        IMAGE_addr <= 1252;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S1269;
      end
      test_b1_S1269: begin
        IMAGE_addr <= 1253;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S1270;
      end
      test_b1_S1270: begin
        IMAGE_addr <= 1254;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S1271;
      end
      test_b1_S1271: begin
        IMAGE_addr <= 1255;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S1272;
      end
      test_b1_S1272: begin
        IMAGE_addr <= 1256;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1273;
      end
      test_b1_S1273: begin
        IMAGE_addr <= 1257;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S1274;
      end
      test_b1_S1274: begin
        IMAGE_addr <= 1258;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S1275;
      end
      test_b1_S1275: begin
        IMAGE_addr <= 1259;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 95;
        test_state <= test_b1_S1276;
      end
      test_b1_S1276: begin
        IMAGE_addr <= 1260;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 95;
        test_state <= test_b1_S1277;
      end
      test_b1_S1277: begin
        IMAGE_addr <= 1261;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 38;
        test_state <= test_b1_S1278;
      end
      test_b1_S1278: begin
        IMAGE_addr <= 1262;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1279;
      end
      test_b1_S1279: begin
        IMAGE_addr <= 1263;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S1280;
      end
      test_b1_S1280: begin
        IMAGE_addr <= 1264;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S1281;
      end
      test_b1_S1281: begin
        IMAGE_addr <= 1265;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S1282;
      end
      test_b1_S1282: begin
        IMAGE_addr <= 1266;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1259;
        test_state <= test_b1_S1283;
      end
      test_b1_S1283: begin
        IMAGE_addr <= 1267;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S1284;
      end
      test_b1_S1284: begin
        IMAGE_addr <= 1268;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S1285;
      end
      test_b1_S1285: begin
        IMAGE_addr <= 1269;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 16;
        test_state <= test_b1_S1286;
      end
      test_b1_S1286: begin
        IMAGE_addr <= 1270;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S1287;
      end
      test_b1_S1287: begin
        IMAGE_addr <= 1271;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 26;
        test_state <= test_b1_S1288;
      end
      test_b1_S1288: begin
        IMAGE_addr <= 1272;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S1289;
      end
      test_b1_S1289: begin
        IMAGE_addr <= 1273;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S1290;
      end
      test_b1_S1290: begin
        IMAGE_addr <= 1274;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S1291;
      end
      test_b1_S1291: begin
        IMAGE_addr <= 1275;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 583;
        test_state <= test_b1_S1292;
      end
      test_b1_S1292: begin
        IMAGE_addr <= 1276;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S1293;
      end
      test_b1_S1293: begin
        IMAGE_addr <= 1277;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S1294;
      end
      test_b1_S1294: begin
        IMAGE_addr <= 1278;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 578;
        test_state <= test_b1_S1295;
      end
      test_b1_S1295: begin
        IMAGE_addr <= 1279;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S1296;
      end
      test_b1_S1296: begin
        IMAGE_addr <= 1280;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S1297;
      end
      test_b1_S1297: begin
        IMAGE_addr <= 1281;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S1298;
      end
      test_b1_S1298: begin
        IMAGE_addr <= 1282;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 400;
        test_state <= test_b1_S1299;
      end
      test_b1_S1299: begin
        IMAGE_addr <= 1283;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1263;
        test_state <= test_b1_S1300;
      end
      test_b1_S1300: begin
        IMAGE_addr <= 1284;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1232;
        test_state <= test_b1_S1301;
      end
      test_b1_S1301: begin
        IMAGE_addr <= 1285;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S1302;
      end
      test_b1_S1302: begin
        IMAGE_addr <= 1286;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1303;
      end
      test_b1_S1303: begin
        IMAGE_addr <= 1287;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 13;
        test_state <= test_b1_S1304;
      end
      test_b1_S1304: begin
        IMAGE_addr <= 1288;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1305;
        test_state <= test_b1_S1305;
      end
      test_b1_S1305: begin
        IMAGE_addr <= 1289;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 583;
        test_state <= test_b1_S1306;
      end
      test_b1_S1306: begin
        IMAGE_addr <= 1290;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S1307;
      end
      test_b1_S1307: begin
        IMAGE_addr <= 1291;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S1308;
      end
      test_b1_S1308: begin
        IMAGE_addr <= 1292;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1259;
        test_state <= test_b1_S1309;
      end
      test_b1_S1309: begin
        IMAGE_addr <= 1293;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1232;
        test_state <= test_b1_S1310;
      end
      test_b1_S1310: begin
        IMAGE_addr <= 1294;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S1311;
      end
      test_b1_S1311: begin
        IMAGE_addr <= 1295;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1312;
      end
      test_b1_S1312: begin
        IMAGE_addr <= 1296;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 13;
        test_state <= test_b1_S1313;
      end
      test_b1_S1313: begin
        IMAGE_addr <= 1297;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1304;
        test_state <= test_b1_S1314;
      end
      test_b1_S1314: begin
        IMAGE_addr <= 1298;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1274;
        test_state <= test_b1_S1315;
      end
      test_b1_S1315: begin
        IMAGE_addr <= 1299;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 286;
        test_state <= test_b1_S1316;
      end
      test_b1_S1316: begin
        IMAGE_addr <= 1300;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S1317;
      end
      test_b1_S1317: begin
        IMAGE_addr <= 1301;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1318;
      end
      test_b1_S1318: begin
        IMAGE_addr <= 1302;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S1319;
      end
      test_b1_S1319: begin
        IMAGE_addr <= 1303;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S1320;
      end
      test_b1_S1320: begin
        IMAGE_addr <= 1304;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S1321;
      end
      test_b1_S1321: begin
        IMAGE_addr <= 1305;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S1322;
      end
      test_b1_S1322: begin
        IMAGE_addr <= 1306;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S1323;
      end
      test_b1_S1323: begin
        IMAGE_addr <= 1307;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4294967295;
        test_state <= test_b1_S1324;
      end
      test_b1_S1324: begin
        IMAGE_addr <= 1308;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S1325;
      end
      test_b1_S1325: begin
        IMAGE_addr <= 1309;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S1326;
      end
      test_b1_S1326: begin
        IMAGE_addr <= 1310;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8;
        test_state <= test_b1_S1327;
      end
      test_b1_S1327: begin
        IMAGE_addr <= 1311;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5734;
        test_state <= test_b1_S1328;
      end
      test_b1_S1328: begin
        IMAGE_addr <= 1312;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 400;
        test_state <= test_b1_S1329;
      end
      test_b1_S1329: begin
        IMAGE_addr <= 1313;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 877;
        test_state <= test_b1_S1330;
      end
      test_b1_S1330: begin
        IMAGE_addr <= 1314;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S1331;
      end
      test_b1_S1331: begin
        IMAGE_addr <= 1315;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S1332;
      end
      test_b1_S1332: begin
        IMAGE_addr <= 1316;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 11;
        test_state <= test_b1_S1333;
      end
      test_b1_S1333: begin
        IMAGE_addr <= 1317;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1319;
        test_state <= test_b1_S1334;
      end
      test_b1_S1334: begin
        IMAGE_addr <= 1318;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1282;
        test_state <= test_b1_S1335;
      end
      test_b1_S1335: begin
        IMAGE_addr <= 1319;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S1336;
      end
      test_b1_S1336: begin
        IMAGE_addr <= 1320;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S1337;
      end
      test_b1_S1337: begin
        IMAGE_addr <= 1321;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1338;
      end
      test_b1_S1338: begin
        IMAGE_addr <= 1322;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1339;
      end
      test_b1_S1339: begin
        IMAGE_addr <= 1323;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1310;
        test_state <= test_b1_S1340;
      end
      test_b1_S1340: begin
        IMAGE_addr <= 1324;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 25;
        test_state <= test_b1_S1341;
      end
      test_b1_S1341: begin
        IMAGE_addr <= 1325;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 52;
        test_state <= test_b1_S1342;
      end
      test_b1_S1342: begin
        IMAGE_addr <= 1326;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 371;
        test_state <= test_b1_S1343;
      end
      test_b1_S1343: begin
        IMAGE_addr <= 1327;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 400;
        test_state <= test_b1_S1344;
      end
      test_b1_S1344: begin
        IMAGE_addr <= 1328;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 391;
        test_state <= test_b1_S1345;
      end
      test_b1_S1345: begin
        IMAGE_addr <= 1329;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S1346;
      end
      test_b1_S1346: begin
        IMAGE_addr <= 1330;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 32;
        test_state <= test_b1_S1347;
      end
      test_b1_S1347: begin
        IMAGE_addr <= 1331;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 359;
        test_state <= test_b1_S1348;
      end
      test_b1_S1348: begin
        IMAGE_addr <= 1332;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S1349;
      end
      test_b1_S1349: begin
        IMAGE_addr <= 1333;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 63;
        test_state <= test_b1_S1350;
      end
      test_b1_S1350: begin
        IMAGE_addr <= 1334;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 359;
        test_state <= test_b1_S1351;
      end
      test_b1_S1351: begin
        IMAGE_addr <= 1335;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 371;
        test_state <= test_b1_S1352;
      end
      test_b1_S1352: begin
        IMAGE_addr <= 1336;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S1353;
      end
      test_b1_S1353: begin
        IMAGE_addr <= 1337;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S1354;
      end
      test_b1_S1354: begin
        IMAGE_addr <= 1338;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1355;
      end
      test_b1_S1355: begin
        IMAGE_addr <= 1339;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1356;
      end
      test_b1_S1356: begin
        IMAGE_addr <= 1340;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S1357;
      end
      test_b1_S1357: begin
        IMAGE_addr <= 1341;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S1358;
      end
      test_b1_S1358: begin
        IMAGE_addr <= 1342;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S1359;
      end
      test_b1_S1359: begin
        IMAGE_addr <= 1343;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 140;
        test_state <= test_b1_S1360;
      end
      test_b1_S1360: begin
        IMAGE_addr <= 1344;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 25;
        test_state <= test_b1_S1361;
      end
      test_b1_S1361: begin
        IMAGE_addr <= 1345;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S1362;
      end
      test_b1_S1362: begin
        IMAGE_addr <= 1346;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 371;
        test_state <= test_b1_S1363;
      end
      test_b1_S1363: begin
        IMAGE_addr <= 1347;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S1364;
      end
      test_b1_S1364: begin
        IMAGE_addr <= 1348;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 29;
        test_state <= test_b1_S1365;
      end
      test_b1_S1365: begin
        IMAGE_addr <= 1349;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 391;
        test_state <= test_b1_S1366;
      end
      test_b1_S1366: begin
        IMAGE_addr <= 1350;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S1367;
      end
      test_b1_S1367: begin
        IMAGE_addr <= 1351;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S1368;
      end
      test_b1_S1368: begin
        IMAGE_addr <= 1352;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1274;
        test_state <= test_b1_S1369;
      end
      test_b1_S1369: begin
        IMAGE_addr <= 1353;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8;
        test_state <= test_b1_S1370;
      end
      test_b1_S1370: begin
        IMAGE_addr <= 1354;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 286;
        test_state <= test_b1_S1371;
      end
      test_b1_S1371: begin
        IMAGE_addr <= 1355;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 400;
        test_state <= test_b1_S1372;
      end
      test_b1_S1372: begin
        IMAGE_addr <= 1356;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1056;
        test_state <= test_b1_S1373;
      end
      test_b1_S1373: begin
        IMAGE_addr <= 1357;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S1374;
      end
      test_b1_S1374: begin
        IMAGE_addr <= 1358;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 310;
        test_state <= test_b1_S1375;
      end
      test_b1_S1375: begin
        IMAGE_addr <= 1359;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 286;
        test_state <= test_b1_S1376;
      end
      test_b1_S1376: begin
        IMAGE_addr <= 1360;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S1377;
      end
      test_b1_S1377: begin
        IMAGE_addr <= 1361;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S1378;
      end
      test_b1_S1378: begin
        IMAGE_addr <= 1362;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 400;
        test_state <= test_b1_S1379;
      end
      test_b1_S1379: begin
        IMAGE_addr <= 1363;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1091;
        test_state <= test_b1_S1380;
      end
      test_b1_S1380: begin
        IMAGE_addr <= 1364;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S1381;
      end
      test_b1_S1381: begin
        IMAGE_addr <= 1365;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1382;
      end
      test_b1_S1382: begin
        IMAGE_addr <= 1366;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 13;
        test_state <= test_b1_S1383;
      end
      test_b1_S1383: begin
        IMAGE_addr <= 1367;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1371;
        test_state <= test_b1_S1384;
      end
      test_b1_S1384: begin
        IMAGE_addr <= 1368;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1355;
        test_state <= test_b1_S1385;
      end
      test_b1_S1385: begin
        IMAGE_addr <= 1369;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S1386;
      end
      test_b1_S1386: begin
        IMAGE_addr <= 1370;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S1387;
      end
      test_b1_S1387: begin
        IMAGE_addr <= 1371;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1321;
        test_state <= test_b1_S1388;
      end
      test_b1_S1388: begin
        IMAGE_addr <= 1372;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S1389;
      end
      test_b1_S1389: begin
        IMAGE_addr <= 1373;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S1390;
      end
      test_b1_S1390: begin
        IMAGE_addr <= 1374;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S1391;
      end
      test_b1_S1391: begin
        IMAGE_addr <= 1375;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1392;
      end
      test_b1_S1392: begin
        IMAGE_addr <= 1376;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 13;
        test_state <= test_b1_S1393;
      end
      test_b1_S1393: begin
        IMAGE_addr <= 1377;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1381;
        test_state <= test_b1_S1394;
      end
      test_b1_S1394: begin
        IMAGE_addr <= 1378;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1352;
        test_state <= test_b1_S1395;
      end
      test_b1_S1395: begin
        IMAGE_addr <= 1379;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S1396;
      end
      test_b1_S1396: begin
        IMAGE_addr <= 1380;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S1397;
      end
      test_b1_S1397: begin
        IMAGE_addr <= 1381;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 52;
        test_state <= test_b1_S1398;
      end
      test_b1_S1398: begin
        IMAGE_addr <= 1382;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1362;
        test_state <= test_b1_S1399;
      end
      test_b1_S1399: begin
        IMAGE_addr <= 1383;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S1400;
      end
      test_b1_S1400: begin
        IMAGE_addr <= 1384;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S1401;
      end
      test_b1_S1401: begin
        IMAGE_addr <= 1385;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1402;
      end
      test_b1_S1402: begin
        IMAGE_addr <= 1386;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1403;
      end
      test_b1_S1403: begin
        IMAGE_addr <= 1387;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1338;
        test_state <= test_b1_S1404;
      end
      test_b1_S1404: begin
        IMAGE_addr <= 1388;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S1405;
      end
      test_b1_S1405: begin
        IMAGE_addr <= 1389;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 32;
        test_state <= test_b1_S1406;
      end
      test_b1_S1406: begin
        IMAGE_addr <= 1390;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 562;
        test_state <= test_b1_S1407;
      end
      test_b1_S1407: begin
        IMAGE_addr <= 1391;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 400;
        test_state <= test_b1_S1408;
      end
      test_b1_S1408: begin
        IMAGE_addr <= 1392;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1232;
        test_state <= test_b1_S1409;
      end
      test_b1_S1409: begin
        IMAGE_addr <= 1393;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1374;
        test_state <= test_b1_S1410;
      end
      test_b1_S1410: begin
        IMAGE_addr <= 1394;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8;
        test_state <= test_b1_S1411;
      end
      test_b1_S1411: begin
        IMAGE_addr <= 1395;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1387;
        test_state <= test_b1_S1412;
      end
      test_b1_S1412: begin
        IMAGE_addr <= 1396;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S1413;
      end
      test_b1_S1413: begin
        IMAGE_addr <= 1397;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S1414;
      end
      test_b1_S1414: begin
        IMAGE_addr <= 1398;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1415;
      end
      test_b1_S1415: begin
        IMAGE_addr <= 1399;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 323;
        test_state <= test_b1_S1416;
      end
      test_b1_S1416: begin
        IMAGE_addr <= 1400;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 37;
        test_state <= test_b1_S1417;
      end
      test_b1_S1417: begin
        IMAGE_addr <= 1401;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 49;
        test_state <= test_b1_S1418;
      end
      test_b1_S1418: begin
        IMAGE_addr <= 1402;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 43;
        test_state <= test_b1_S1419;
      end
      test_b1_S1419: begin
        IMAGE_addr <= 1403;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1420;
      end
      test_b1_S1420: begin
        IMAGE_addr <= 1404;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1398;
        test_state <= test_b1_S1421;
      end
      test_b1_S1421: begin
        IMAGE_addr <= 1405;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 323;
        test_state <= test_b1_S1422;
      end
      test_b1_S1422: begin
        IMAGE_addr <= 1406;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 42;
        test_state <= test_b1_S1423;
      end
      test_b1_S1423: begin
        IMAGE_addr <= 1407;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 49;
        test_state <= test_b1_S1424;
      end
      test_b1_S1424: begin
        IMAGE_addr <= 1408;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 45;
        test_state <= test_b1_S1425;
      end
      test_b1_S1425: begin
        IMAGE_addr <= 1409;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1426;
      end
      test_b1_S1426: begin
        IMAGE_addr <= 1410;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1404;
        test_state <= test_b1_S1427;
      end
      test_b1_S1427: begin
        IMAGE_addr <= 1411;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 323;
        test_state <= test_b1_S1428;
      end
      test_b1_S1428: begin
        IMAGE_addr <= 1412;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 47;
        test_state <= test_b1_S1429;
      end
      test_b1_S1429: begin
        IMAGE_addr <= 1413;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S1430;
      end
      test_b1_S1430: begin
        IMAGE_addr <= 1414;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 119;
        test_state <= test_b1_S1431;
      end
      test_b1_S1431: begin
        IMAGE_addr <= 1415;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S1432;
      end
      test_b1_S1432: begin
        IMAGE_addr <= 1416;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 112;
        test_state <= test_b1_S1433;
      end
      test_b1_S1433: begin
        IMAGE_addr <= 1417;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1434;
      end
      test_b1_S1434: begin
        IMAGE_addr <= 1418;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1410;
        test_state <= test_b1_S1435;
      end
      test_b1_S1435: begin
        IMAGE_addr <= 1419;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 323;
        test_state <= test_b1_S1436;
      end
      test_b1_S1436: begin
        IMAGE_addr <= 1420;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 52;
        test_state <= test_b1_S1437;
      end
      test_b1_S1437: begin
        IMAGE_addr <= 1421;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 100;
        test_state <= test_b1_S1438;
      end
      test_b1_S1438: begin
        IMAGE_addr <= 1422;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S1439;
      end
      test_b1_S1439: begin
        IMAGE_addr <= 1423;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 111;
        test_state <= test_b1_S1440;
      end
      test_b1_S1440: begin
        IMAGE_addr <= 1424;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 112;
        test_state <= test_b1_S1441;
      end
      test_b1_S1441: begin
        IMAGE_addr <= 1425;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1442;
      end
      test_b1_S1442: begin
        IMAGE_addr <= 1426;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1418;
        test_state <= test_b1_S1443;
      end
      test_b1_S1443: begin
        IMAGE_addr <= 1427;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 323;
        test_state <= test_b1_S1444;
      end
      test_b1_S1444: begin
        IMAGE_addr <= 1428;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 57;
        test_state <= test_b1_S1445;
      end
      test_b1_S1445: begin
        IMAGE_addr <= 1429;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S1446;
      end
      test_b1_S1446: begin
        IMAGE_addr <= 1430;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 110;
        test_state <= test_b1_S1447;
      end
      test_b1_S1447: begin
        IMAGE_addr <= 1431;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 100;
        test_state <= test_b1_S1448;
      end
      test_b1_S1448: begin
        IMAGE_addr <= 1432;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1449;
      end
      test_b1_S1449: begin
        IMAGE_addr <= 1433;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1426;
        test_state <= test_b1_S1450;
      end
      test_b1_S1450: begin
        IMAGE_addr <= 1434;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 323;
        test_state <= test_b1_S1451;
      end
      test_b1_S1451: begin
        IMAGE_addr <= 1435;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 62;
        test_state <= test_b1_S1452;
      end
      test_b1_S1452: begin
        IMAGE_addr <= 1436;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 111;
        test_state <= test_b1_S1453;
      end
      test_b1_S1453: begin
        IMAGE_addr <= 1437;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S1454;
      end
      test_b1_S1454: begin
        IMAGE_addr <= 1438;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1455;
      end
      test_b1_S1455: begin
        IMAGE_addr <= 1439;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1433;
        test_state <= test_b1_S1456;
      end
      test_b1_S1456: begin
        IMAGE_addr <= 1440;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 323;
        test_state <= test_b1_S1457;
      end
      test_b1_S1457: begin
        IMAGE_addr <= 1441;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 67;
        test_state <= test_b1_S1458;
      end
      test_b1_S1458: begin
        IMAGE_addr <= 1442;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 120;
        test_state <= test_b1_S1459;
      end
      test_b1_S1459: begin
        IMAGE_addr <= 1443;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 111;
        test_state <= test_b1_S1460;
      end
      test_b1_S1460: begin
        IMAGE_addr <= 1444;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S1461;
      end
      test_b1_S1461: begin
        IMAGE_addr <= 1445;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1462;
      end
      test_b1_S1462: begin
        IMAGE_addr <= 1446;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1439;
        test_state <= test_b1_S1463;
      end
      test_b1_S1463: begin
        IMAGE_addr <= 1447;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 323;
        test_state <= test_b1_S1464;
      end
      test_b1_S1464: begin
        IMAGE_addr <= 1448;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 72;
        test_state <= test_b1_S1465;
      end
      test_b1_S1465: begin
        IMAGE_addr <= 1449;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 64;
        test_state <= test_b1_S1466;
      end
      test_b1_S1466: begin
        IMAGE_addr <= 1450;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1467;
      end
      test_b1_S1467: begin
        IMAGE_addr <= 1451;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1446;
        test_state <= test_b1_S1468;
      end
      test_b1_S1468: begin
        IMAGE_addr <= 1452;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 323;
        test_state <= test_b1_S1469;
      end
      test_b1_S1469: begin
        IMAGE_addr <= 1453;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 77;
        test_state <= test_b1_S1470;
      end
      test_b1_S1470: begin
        IMAGE_addr <= 1454;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 33;
        test_state <= test_b1_S1471;
      end
      test_b1_S1471: begin
        IMAGE_addr <= 1455;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1472;
      end
      test_b1_S1472: begin
        IMAGE_addr <= 1456;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1451;
        test_state <= test_b1_S1473;
      end
      test_b1_S1473: begin
        IMAGE_addr <= 1457;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 323;
        test_state <= test_b1_S1474;
      end
      test_b1_S1474: begin
        IMAGE_addr <= 1458;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 82;
        test_state <= test_b1_S1475;
      end
      test_b1_S1475: begin
        IMAGE_addr <= 1459;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 43;
        test_state <= test_b1_S1476;
      end
      test_b1_S1476: begin
        IMAGE_addr <= 1460;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1477;
      end
      test_b1_S1477: begin
        IMAGE_addr <= 1461;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1456;
        test_state <= test_b1_S1478;
      end
      test_b1_S1478: begin
        IMAGE_addr <= 1462;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 323;
        test_state <= test_b1_S1479;
      end
      test_b1_S1479: begin
        IMAGE_addr <= 1463;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 87;
        test_state <= test_b1_S1480;
      end
      test_b1_S1480: begin
        IMAGE_addr <= 1464;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 45;
        test_state <= test_b1_S1481;
      end
      test_b1_S1481: begin
        IMAGE_addr <= 1465;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1482;
      end
      test_b1_S1482: begin
        IMAGE_addr <= 1466;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1461;
        test_state <= test_b1_S1483;
      end
      test_b1_S1483: begin
        IMAGE_addr <= 1467;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 323;
        test_state <= test_b1_S1484;
      end
      test_b1_S1484: begin
        IMAGE_addr <= 1468;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 92;
        test_state <= test_b1_S1485;
      end
      test_b1_S1485: begin
        IMAGE_addr <= 1469;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 42;
        test_state <= test_b1_S1486;
      end
      test_b1_S1486: begin
        IMAGE_addr <= 1470;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1487;
      end
      test_b1_S1487: begin
        IMAGE_addr <= 1471;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1466;
        test_state <= test_b1_S1488;
      end
      test_b1_S1488: begin
        IMAGE_addr <= 1472;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 323;
        test_state <= test_b1_S1489;
      end
      test_b1_S1489: begin
        IMAGE_addr <= 1473;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S1490;
      end
      test_b1_S1490: begin
        IMAGE_addr <= 1474;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 47;
        test_state <= test_b1_S1491;
      end
      test_b1_S1491: begin
        IMAGE_addr <= 1475;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 109;
        test_state <= test_b1_S1492;
      end
      test_b1_S1492: begin
        IMAGE_addr <= 1476;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 111;
        test_state <= test_b1_S1493;
      end
      test_b1_S1493: begin
        IMAGE_addr <= 1477;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 100;
        test_state <= test_b1_S1494;
      end
      test_b1_S1494: begin
        IMAGE_addr <= 1478;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1495;
      end
      test_b1_S1495: begin
        IMAGE_addr <= 1479;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1471;
        test_state <= test_b1_S1496;
      end
      test_b1_S1496: begin
        IMAGE_addr <= 1480;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 323;
        test_state <= test_b1_S1497;
      end
      test_b1_S1497: begin
        IMAGE_addr <= 1481;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 102;
        test_state <= test_b1_S1498;
      end
      test_b1_S1498: begin
        IMAGE_addr <= 1482;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 60;
        test_state <= test_b1_S1499;
      end
      test_b1_S1499: begin
        IMAGE_addr <= 1483;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 60;
        test_state <= test_b1_S1500;
      end
      test_b1_S1500: begin
        IMAGE_addr <= 1484;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1501;
      end
      test_b1_S1501: begin
        IMAGE_addr <= 1485;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1479;
        test_state <= test_b1_S1502;
      end
      test_b1_S1502: begin
        IMAGE_addr <= 1486;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 323;
        test_state <= test_b1_S1503;
      end
      test_b1_S1503: begin
        IMAGE_addr <= 1487;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 107;
        test_state <= test_b1_S1504;
      end
      test_b1_S1504: begin
        IMAGE_addr <= 1488;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 62;
        test_state <= test_b1_S1505;
      end
      test_b1_S1505: begin
        IMAGE_addr <= 1489;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 62;
        test_state <= test_b1_S1506;
      end
      test_b1_S1506: begin
        IMAGE_addr <= 1490;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1507;
      end
      test_b1_S1507: begin
        IMAGE_addr <= 1491;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1485;
        test_state <= test_b1_S1508;
      end
      test_b1_S1508: begin
        IMAGE_addr <= 1492;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S1509;
      end
      test_b1_S1509: begin
        IMAGE_addr <= 1493;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 400;
        test_state <= test_b1_S1510;
      end
      test_b1_S1510: begin
        IMAGE_addr <= 1494;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S1511;
      end
      test_b1_S1511: begin
        IMAGE_addr <= 1495;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S1512;
      end
      test_b1_S1512: begin
        IMAGE_addr <= 1496;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 98;
        test_state <= test_b1_S1513;
      end
      test_b1_S1513: begin
        IMAGE_addr <= 1497;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1514;
      end
      test_b1_S1514: begin
        IMAGE_addr <= 1498;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1491;
        test_state <= test_b1_S1515;
      end
      test_b1_S1515: begin
        IMAGE_addr <= 1499;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 323;
        test_state <= test_b1_S1516;
      end
      test_b1_S1516: begin
        IMAGE_addr <= 1500;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 32;
        test_state <= test_b1_S1517;
      end
      test_b1_S1517: begin
        IMAGE_addr <= 1501;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 100;
        test_state <= test_b1_S1518;
      end
      test_b1_S1518: begin
        IMAGE_addr <= 1502;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 117;
        test_state <= test_b1_S1519;
      end
      test_b1_S1519: begin
        IMAGE_addr <= 1503;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 112;
        test_state <= test_b1_S1520;
      end
      test_b1_S1520: begin
        IMAGE_addr <= 1504;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1521;
      end
      test_b1_S1521: begin
        IMAGE_addr <= 1505;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1498;
        test_state <= test_b1_S1522;
      end
      test_b1_S1522: begin
        IMAGE_addr <= 1506;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 323;
        test_state <= test_b1_S1523;
      end
      test_b1_S1523: begin
        IMAGE_addr <= 1507;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 117;
        test_state <= test_b1_S1524;
      end
      test_b1_S1524: begin
        IMAGE_addr <= 1508;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S1525;
      end
      test_b1_S1525: begin
        IMAGE_addr <= 1509;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 110;
        test_state <= test_b1_S1526;
      end
      test_b1_S1526: begin
        IMAGE_addr <= 1510;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1527;
      end
      test_b1_S1527: begin
        IMAGE_addr <= 1511;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1505;
        test_state <= test_b1_S1528;
      end
      test_b1_S1528: begin
        IMAGE_addr <= 1512;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 323;
        test_state <= test_b1_S1529;
      end
      test_b1_S1529: begin
        IMAGE_addr <= 1513;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 112;
        test_state <= test_b1_S1530;
      end
      test_b1_S1530: begin
        IMAGE_addr <= 1514;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 111;
        test_state <= test_b1_S1531;
      end
      test_b1_S1531: begin
        IMAGE_addr <= 1515;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 117;
        test_state <= test_b1_S1532;
      end
      test_b1_S1532: begin
        IMAGE_addr <= 1516;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S1533;
      end
      test_b1_S1533: begin
        IMAGE_addr <= 1517;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1534;
      end
      test_b1_S1534: begin
        IMAGE_addr <= 1518;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1511;
        test_state <= test_b1_S1535;
      end
      test_b1_S1535: begin
        IMAGE_addr <= 1519;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S1536;
      end
      test_b1_S1536: begin
        IMAGE_addr <= 1520;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 562;
        test_state <= test_b1_S1537;
      end
      test_b1_S1537: begin
        IMAGE_addr <= 1521;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S1538;
      end
      test_b1_S1538: begin
        IMAGE_addr <= 1522;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 99;
        test_state <= test_b1_S1539;
      end
      test_b1_S1539: begin
        IMAGE_addr <= 1523;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 99;
        test_state <= test_b1_S1540;
      end
      test_b1_S1540: begin
        IMAGE_addr <= 1524;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S1541;
      end
      test_b1_S1541: begin
        IMAGE_addr <= 1525;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 112;
        test_state <= test_b1_S1542;
      end
      test_b1_S1542: begin
        IMAGE_addr <= 1526;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S1543;
      end
      test_b1_S1543: begin
        IMAGE_addr <= 1527;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1544;
      end
      test_b1_S1544: begin
        IMAGE_addr <= 1528;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1518;
        test_state <= test_b1_S1545;
      end
      test_b1_S1545: begin
        IMAGE_addr <= 1529;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S1546;
      end
      test_b1_S1546: begin
        IMAGE_addr <= 1530;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 206;
        test_state <= test_b1_S1547;
      end
      test_b1_S1547: begin
        IMAGE_addr <= 1531;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 104;
        test_state <= test_b1_S1548;
      end
      test_b1_S1548: begin
        IMAGE_addr <= 1532;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S1549;
      end
      test_b1_S1549: begin
        IMAGE_addr <= 1533;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S1550;
      end
      test_b1_S1550: begin
        IMAGE_addr <= 1534;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S1551;
      end
      test_b1_S1551: begin
        IMAGE_addr <= 1535;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1552;
      end
      test_b1_S1552: begin
        IMAGE_addr <= 1536;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1528;
        test_state <= test_b1_S1553;
      end
      test_b1_S1553: begin
        IMAGE_addr <= 1537;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S1554;
      end
      test_b1_S1554: begin
        IMAGE_addr <= 1538;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 213;
        test_state <= test_b1_S1555;
      end
      test_b1_S1555: begin
        IMAGE_addr <= 1539;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 44;
        test_state <= test_b1_S1556;
      end
      test_b1_S1556: begin
        IMAGE_addr <= 1540;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1557;
      end
      test_b1_S1557: begin
        IMAGE_addr <= 1541;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1536;
        test_state <= test_b1_S1558;
      end
      test_b1_S1558: begin
        IMAGE_addr <= 1542;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S1559;
      end
      test_b1_S1559: begin
        IMAGE_addr <= 1543;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 621;
        test_state <= test_b1_S1560;
      end
      test_b1_S1560: begin
        IMAGE_addr <= 1544;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 99;
        test_state <= test_b1_S1561;
      end
      test_b1_S1561: begin
        IMAGE_addr <= 1545;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S1562;
      end
      test_b1_S1562: begin
        IMAGE_addr <= 1546;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S1563;
      end
      test_b1_S1563: begin
        IMAGE_addr <= 1547;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S1564;
      end
      test_b1_S1564: begin
        IMAGE_addr <= 1548;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S1565;
      end
      test_b1_S1565: begin
        IMAGE_addr <= 1549;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S1566;
      end
      test_b1_S1566: begin
        IMAGE_addr <= 1550;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1567;
      end
      test_b1_S1567: begin
        IMAGE_addr <= 1551;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1541;
        test_state <= test_b1_S1568;
      end
      test_b1_S1568: begin
        IMAGE_addr <= 1552;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S1569;
      end
      test_b1_S1569: begin
        IMAGE_addr <= 1553;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 637;
        test_state <= test_b1_S1570;
      end
      test_b1_S1570: begin
        IMAGE_addr <= 1554;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 93;
        test_state <= test_b1_S1571;
      end
      test_b1_S1571: begin
        IMAGE_addr <= 1555;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 93;
        test_state <= test_b1_S1572;
      end
      test_b1_S1572: begin
        IMAGE_addr <= 1556;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1573;
      end
      test_b1_S1573: begin
        IMAGE_addr <= 1557;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1551;
        test_state <= test_b1_S1574;
      end
      test_b1_S1574: begin
        IMAGE_addr <= 1558;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S1575;
      end
      test_b1_S1575: begin
        IMAGE_addr <= 1559;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 659;
        test_state <= test_b1_S1576;
      end
      test_b1_S1576: begin
        IMAGE_addr <= 1560;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 58;
        test_state <= test_b1_S1577;
      end
      test_b1_S1577: begin
        IMAGE_addr <= 1561;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1578;
      end
      test_b1_S1578: begin
        IMAGE_addr <= 1562;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1557;
        test_state <= test_b1_S1579;
      end
      test_b1_S1579: begin
        IMAGE_addr <= 1563;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S1580;
      end
      test_b1_S1580: begin
        IMAGE_addr <= 1564;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 596;
        test_state <= test_b1_S1581;
      end
      test_b1_S1581: begin
        IMAGE_addr <= 1565;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 104;
        test_state <= test_b1_S1582;
      end
      test_b1_S1582: begin
        IMAGE_addr <= 1566;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S1583;
      end
      test_b1_S1583: begin
        IMAGE_addr <= 1567;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S1584;
      end
      test_b1_S1584: begin
        IMAGE_addr <= 1568;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 100;
        test_state <= test_b1_S1585;
      end
      test_b1_S1585: begin
        IMAGE_addr <= 1569;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S1586;
      end
      test_b1_S1586: begin
        IMAGE_addr <= 1570;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S1587;
      end
      test_b1_S1587: begin
        IMAGE_addr <= 1571;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1588;
      end
      test_b1_S1588: begin
        IMAGE_addr <= 1572;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1562;
        test_state <= test_b1_S1589;
      end
      test_b1_S1589: begin
        IMAGE_addr <= 1573;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S1590;
      end
      test_b1_S1590: begin
        IMAGE_addr <= 1574;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 371;
        test_state <= test_b1_S1591;
      end
      test_b1_S1591: begin
        IMAGE_addr <= 1575;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 99;
        test_state <= test_b1_S1592;
      end
      test_b1_S1592: begin
        IMAGE_addr <= 1576;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S1593;
      end
      test_b1_S1593: begin
        IMAGE_addr <= 1577;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1594;
      end
      test_b1_S1594: begin
        IMAGE_addr <= 1578;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1572;
        test_state <= test_b1_S1595;
      end
      test_b1_S1595: begin
        IMAGE_addr <= 1579;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S1596;
      end
      test_b1_S1596: begin
        IMAGE_addr <= 1580;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 359;
        test_state <= test_b1_S1597;
      end
      test_b1_S1597: begin
        IMAGE_addr <= 1581;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 112;
        test_state <= test_b1_S1598;
      end
      test_b1_S1598: begin
        IMAGE_addr <= 1582;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 117;
        test_state <= test_b1_S1599;
      end
      test_b1_S1599: begin
        IMAGE_addr <= 1583;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S1600;
      end
      test_b1_S1600: begin
        IMAGE_addr <= 1584;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 99;
        test_state <= test_b1_S1601;
      end
      test_b1_S1601: begin
        IMAGE_addr <= 1585;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1602;
      end
      test_b1_S1602: begin
        IMAGE_addr <= 1586;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1578;
        test_state <= test_b1_S1603;
      end
      test_b1_S1603: begin
        IMAGE_addr <= 1587;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S1604;
      end
      test_b1_S1604: begin
        IMAGE_addr <= 1588;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 407;
        test_state <= test_b1_S1605;
      end
      test_b1_S1605: begin
        IMAGE_addr <= 1589;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S1606;
      end
      test_b1_S1606: begin
        IMAGE_addr <= 1590;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S1607;
      end
      test_b1_S1607: begin
        IMAGE_addr <= 1591;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 109;
        test_state <= test_b1_S1608;
      end
      test_b1_S1608: begin
        IMAGE_addr <= 1592;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S1609;
      end
      test_b1_S1609: begin
        IMAGE_addr <= 1593;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 112;
        test_state <= test_b1_S1610;
      end
      test_b1_S1610: begin
        IMAGE_addr <= 1594;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 75;
        test_state <= test_b1_S1611;
      end
      test_b1_S1611: begin
        IMAGE_addr <= 1595;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S1612;
      end
      test_b1_S1612: begin
        IMAGE_addr <= 1596;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 121;
        test_state <= test_b1_S1613;
      end
      test_b1_S1613: begin
        IMAGE_addr <= 1597;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S1614;
      end
      test_b1_S1614: begin
        IMAGE_addr <= 1598;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1615;
      end
      test_b1_S1615: begin
        IMAGE_addr <= 1599;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1586;
        test_state <= test_b1_S1616;
      end
      test_b1_S1616: begin
        IMAGE_addr <= 1600;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S1617;
      end
      test_b1_S1617: begin
        IMAGE_addr <= 1601;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 385;
        test_state <= test_b1_S1618;
      end
      test_b1_S1618: begin
        IMAGE_addr <= 1602;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 60;
        test_state <= test_b1_S1619;
      end
      test_b1_S1619: begin
        IMAGE_addr <= 1603;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 112;
        test_state <= test_b1_S1620;
      end
      test_b1_S1620: begin
        IMAGE_addr <= 1604;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 117;
        test_state <= test_b1_S1621;
      end
      test_b1_S1621: begin
        IMAGE_addr <= 1605;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S1622;
      end
      test_b1_S1622: begin
        IMAGE_addr <= 1606;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S1623;
      end
      test_b1_S1623: begin
        IMAGE_addr <= 1607;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 62;
        test_state <= test_b1_S1624;
      end
      test_b1_S1624: begin
        IMAGE_addr <= 1608;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1625;
      end
      test_b1_S1625: begin
        IMAGE_addr <= 1609;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1599;
        test_state <= test_b1_S1626;
      end
      test_b1_S1626: begin
        IMAGE_addr <= 1610;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S1627;
      end
      test_b1_S1627: begin
        IMAGE_addr <= 1611;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 132;
        test_state <= test_b1_S1628;
      end
      test_b1_S1628: begin
        IMAGE_addr <= 1612;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 111;
        test_state <= test_b1_S1629;
      end
      test_b1_S1629: begin
        IMAGE_addr <= 1613;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 118;
        test_state <= test_b1_S1630;
      end
      test_b1_S1630: begin
        IMAGE_addr <= 1614;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S1631;
      end
      test_b1_S1631: begin
        IMAGE_addr <= 1615;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S1632;
      end
      test_b1_S1632: begin
        IMAGE_addr <= 1616;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1633;
      end
      test_b1_S1633: begin
        IMAGE_addr <= 1617;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1609;
        test_state <= test_b1_S1634;
      end
      test_b1_S1634: begin
        IMAGE_addr <= 1618;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S1635;
      end
      test_b1_S1635: begin
        IMAGE_addr <= 1619;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S1636;
      end
      test_b1_S1636: begin
        IMAGE_addr <= 1620;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 113;
        test_state <= test_b1_S1637;
      end
      test_b1_S1637: begin
        IMAGE_addr <= 1621;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 117;
        test_state <= test_b1_S1638;
      end
      test_b1_S1638: begin
        IMAGE_addr <= 1622;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 111;
        test_state <= test_b1_S1639;
      end
      test_b1_S1639: begin
        IMAGE_addr <= 1623;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S1640;
      end
      test_b1_S1640: begin
        IMAGE_addr <= 1624;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S1641;
      end
      test_b1_S1641: begin
        IMAGE_addr <= 1625;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1642;
      end
      test_b1_S1642: begin
        IMAGE_addr <= 1626;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1617;
        test_state <= test_b1_S1643;
      end
      test_b1_S1643: begin
        IMAGE_addr <= 1627;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S1644;
      end
      test_b1_S1644: begin
        IMAGE_addr <= 1628;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 140;
        test_state <= test_b1_S1645;
      end
      test_b1_S1645: begin
        IMAGE_addr <= 1629;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 110;
        test_state <= test_b1_S1646;
      end
      test_b1_S1646: begin
        IMAGE_addr <= 1630;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 111;
        test_state <= test_b1_S1647;
      end
      test_b1_S1647: begin
        IMAGE_addr <= 1631;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S1648;
      end
      test_b1_S1648: begin
        IMAGE_addr <= 1632;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1649;
      end
      test_b1_S1649: begin
        IMAGE_addr <= 1633;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1626;
        test_state <= test_b1_S1650;
      end
      test_b1_S1650: begin
        IMAGE_addr <= 1634;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S1651;
      end
      test_b1_S1651: begin
        IMAGE_addr <= 1635;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 147;
        test_state <= test_b1_S1652;
      end
      test_b1_S1652: begin
        IMAGE_addr <= 1636;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 111;
        test_state <= test_b1_S1653;
      end
      test_b1_S1653: begin
        IMAGE_addr <= 1637;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 110;
        test_state <= test_b1_S1654;
      end
      test_b1_S1654: begin
        IMAGE_addr <= 1638;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1655;
      end
      test_b1_S1655: begin
        IMAGE_addr <= 1639;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1633;
        test_state <= test_b1_S1656;
      end
      test_b1_S1656: begin
        IMAGE_addr <= 1640;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S1657;
      end
      test_b1_S1657: begin
        IMAGE_addr <= 1641;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 155;
        test_state <= test_b1_S1658;
      end
      test_b1_S1658: begin
        IMAGE_addr <= 1642;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 111;
        test_state <= test_b1_S1659;
      end
      test_b1_S1659: begin
        IMAGE_addr <= 1643;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 102;
        test_state <= test_b1_S1660;
      end
      test_b1_S1660: begin
        IMAGE_addr <= 1644;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 102;
        test_state <= test_b1_S1661;
      end
      test_b1_S1661: begin
        IMAGE_addr <= 1645;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1662;
      end
      test_b1_S1662: begin
        IMAGE_addr <= 1646;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1639;
        test_state <= test_b1_S1663;
      end
      test_b1_S1663: begin
        IMAGE_addr <= 1647;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S1664;
      end
      test_b1_S1664: begin
        IMAGE_addr <= 1648;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 163;
        test_state <= test_b1_S1665;
      end
      test_b1_S1665: begin
        IMAGE_addr <= 1649;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 47;
        test_state <= test_b1_S1666;
      end
      test_b1_S1666: begin
        IMAGE_addr <= 1650;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1667;
      end
      test_b1_S1667: begin
        IMAGE_addr <= 1651;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1646;
        test_state <= test_b1_S1668;
      end
      test_b1_S1668: begin
        IMAGE_addr <= 1652;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S1669;
      end
      test_b1_S1669: begin
        IMAGE_addr <= 1653;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 170;
        test_state <= test_b1_S1670;
      end
      test_b1_S1670: begin
        IMAGE_addr <= 1654;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 109;
        test_state <= test_b1_S1671;
      end
      test_b1_S1671: begin
        IMAGE_addr <= 1655;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 111;
        test_state <= test_b1_S1672;
      end
      test_b1_S1672: begin
        IMAGE_addr <= 1656;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 100;
        test_state <= test_b1_S1673;
      end
      test_b1_S1673: begin
        IMAGE_addr <= 1657;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1674;
      end
      test_b1_S1674: begin
        IMAGE_addr <= 1658;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1651;
        test_state <= test_b1_S1675;
      end
      test_b1_S1675: begin
        IMAGE_addr <= 1659;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S1676;
      end
      test_b1_S1676: begin
        IMAGE_addr <= 1660;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 176;
        test_state <= test_b1_S1677;
      end
      test_b1_S1677: begin
        IMAGE_addr <= 1661;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 110;
        test_state <= test_b1_S1678;
      end
      test_b1_S1678: begin
        IMAGE_addr <= 1662;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S1679;
      end
      test_b1_S1679: begin
        IMAGE_addr <= 1663;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 103;
        test_state <= test_b1_S1680;
      end
      test_b1_S1680: begin
        IMAGE_addr <= 1664;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S1681;
      end
      test_b1_S1681: begin
        IMAGE_addr <= 1665;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S1682;
      end
      test_b1_S1682: begin
        IMAGE_addr <= 1666;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S1683;
      end
      test_b1_S1683: begin
        IMAGE_addr <= 1667;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1684;
      end
      test_b1_S1684: begin
        IMAGE_addr <= 1668;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1658;
        test_state <= test_b1_S1685;
      end
      test_b1_S1685: begin
        IMAGE_addr <= 1669;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S1686;
      end
      test_b1_S1686: begin
        IMAGE_addr <= 1670;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 183;
        test_state <= test_b1_S1687;
      end
      test_b1_S1687: begin
        IMAGE_addr <= 1671;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 100;
        test_state <= test_b1_S1688;
      end
      test_b1_S1688: begin
        IMAGE_addr <= 1672;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 111;
        test_state <= test_b1_S1689;
      end
      test_b1_S1689: begin
        IMAGE_addr <= 1673;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1690;
      end
      test_b1_S1690: begin
        IMAGE_addr <= 1674;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1668;
        test_state <= test_b1_S1691;
      end
      test_b1_S1691: begin
        IMAGE_addr <= 1675;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S1692;
      end
      test_b1_S1692: begin
        IMAGE_addr <= 1676;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 943;
        test_state <= test_b1_S1693;
      end
      test_b1_S1693: begin
        IMAGE_addr <= 1677;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 110;
        test_state <= test_b1_S1694;
      end
      test_b1_S1694: begin
        IMAGE_addr <= 1678;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 117;
        test_state <= test_b1_S1695;
      end
      test_b1_S1695: begin
        IMAGE_addr <= 1679;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 109;
        test_state <= test_b1_S1696;
      end
      test_b1_S1696: begin
        IMAGE_addr <= 1680;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 98;
        test_state <= test_b1_S1697;
      end
      test_b1_S1697: begin
        IMAGE_addr <= 1681;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S1698;
      end
      test_b1_S1698: begin
        IMAGE_addr <= 1682;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S1699;
      end
      test_b1_S1699: begin
        IMAGE_addr <= 1683;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S1700;
      end
      test_b1_S1700: begin
        IMAGE_addr <= 1684;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1701;
      end
      test_b1_S1701: begin
        IMAGE_addr <= 1685;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1674;
        test_state <= test_b1_S1702;
      end
      test_b1_S1702: begin
        IMAGE_addr <= 1686;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S1703;
      end
      test_b1_S1703: begin
        IMAGE_addr <= 1687;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 122;
        test_state <= test_b1_S1704;
      end
      test_b1_S1704: begin
        IMAGE_addr <= 1688;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 119;
        test_state <= test_b1_S1705;
      end
      test_b1_S1705: begin
        IMAGE_addr <= 1689;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S1706;
      end
      test_b1_S1706: begin
        IMAGE_addr <= 1690;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S1707;
      end
      test_b1_S1707: begin
        IMAGE_addr <= 1691;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S1708;
      end
      test_b1_S1708: begin
        IMAGE_addr <= 1692;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1709;
      end
      test_b1_S1709: begin
        IMAGE_addr <= 1693;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1685;
        test_state <= test_b1_S1710;
      end
      test_b1_S1710: begin
        IMAGE_addr <= 1694;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S1711;
      end
      test_b1_S1711: begin
        IMAGE_addr <= 1695;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1239;
        test_state <= test_b1_S1712;
      end
      test_b1_S1712: begin
        IMAGE_addr <= 1696;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 39;
        test_state <= test_b1_S1713;
      end
      test_b1_S1713: begin
        IMAGE_addr <= 1697;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1714;
      end
      test_b1_S1714: begin
        IMAGE_addr <= 1698;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1693;
        test_state <= test_b1_S1715;
      end
      test_b1_S1715: begin
        IMAGE_addr <= 1699;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S1716;
      end
      test_b1_S1716: begin
        IMAGE_addr <= 1700;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 189;
        test_state <= test_b1_S1717;
      end
      test_b1_S1717: begin
        IMAGE_addr <= 1701;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 64;
        test_state <= test_b1_S1718;
      end
      test_b1_S1718: begin
        IMAGE_addr <= 1702;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 43;
        test_state <= test_b1_S1719;
      end
      test_b1_S1719: begin
        IMAGE_addr <= 1703;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1720;
      end
      test_b1_S1720: begin
        IMAGE_addr <= 1704;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1698;
        test_state <= test_b1_S1721;
      end
      test_b1_S1721: begin
        IMAGE_addr <= 1705;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S1722;
      end
      test_b1_S1722: begin
        IMAGE_addr <= 1706;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 197;
        test_state <= test_b1_S1723;
      end
      test_b1_S1723: begin
        IMAGE_addr <= 1707;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 33;
        test_state <= test_b1_S1724;
      end
      test_b1_S1724: begin
        IMAGE_addr <= 1708;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 43;
        test_state <= test_b1_S1725;
      end
      test_b1_S1725: begin
        IMAGE_addr <= 1709;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1726;
      end
      test_b1_S1726: begin
        IMAGE_addr <= 1710;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1704;
        test_state <= test_b1_S1727;
      end
      test_b1_S1727: begin
        IMAGE_addr <= 1711;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S1728;
      end
      test_b1_S1728: begin
        IMAGE_addr <= 1712;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 892;
        test_state <= test_b1_S1729;
      end
      test_b1_S1729: begin
        IMAGE_addr <= 1713;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 107;
        test_state <= test_b1_S1730;
      end
      test_b1_S1730: begin
        IMAGE_addr <= 1714;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S1731;
      end
      test_b1_S1731: begin
        IMAGE_addr <= 1715;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S1732;
      end
      test_b1_S1732: begin
        IMAGE_addr <= 1716;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 112;
        test_state <= test_b1_S1733;
      end
      test_b1_S1733: begin
        IMAGE_addr <= 1717;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 83;
        test_state <= test_b1_S1734;
      end
      test_b1_S1734: begin
        IMAGE_addr <= 1718;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S1735;
      end
      test_b1_S1735: begin
        IMAGE_addr <= 1719;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S1736;
      end
      test_b1_S1736: begin
        IMAGE_addr <= 1720;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S1737;
      end
      test_b1_S1737: begin
        IMAGE_addr <= 1721;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 110;
        test_state <= test_b1_S1738;
      end
      test_b1_S1738: begin
        IMAGE_addr <= 1722;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 103;
        test_state <= test_b1_S1739;
      end
      test_b1_S1739: begin
        IMAGE_addr <= 1723;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1740;
      end
      test_b1_S1740: begin
        IMAGE_addr <= 1724;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1710;
        test_state <= test_b1_S1741;
      end
      test_b1_S1741: begin
        IMAGE_addr <= 1725;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S1742;
      end
      test_b1_S1742: begin
        IMAGE_addr <= 1726;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 877;
        test_state <= test_b1_S1743;
      end
      test_b1_S1743: begin
        IMAGE_addr <= 1727;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 103;
        test_state <= test_b1_S1744;
      end
      test_b1_S1744: begin
        IMAGE_addr <= 1728;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S1745;
      end
      test_b1_S1745: begin
        IMAGE_addr <= 1729;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S1746;
      end
      test_b1_S1746: begin
        IMAGE_addr <= 1730;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 76;
        test_state <= test_b1_S1747;
      end
      test_b1_S1747: begin
        IMAGE_addr <= 1731;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S1748;
      end
      test_b1_S1748: begin
        IMAGE_addr <= 1732;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 110;
        test_state <= test_b1_S1749;
      end
      test_b1_S1749: begin
        IMAGE_addr <= 1733;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 103;
        test_state <= test_b1_S1750;
      end
      test_b1_S1750: begin
        IMAGE_addr <= 1734;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S1751;
      end
      test_b1_S1751: begin
        IMAGE_addr <= 1735;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 104;
        test_state <= test_b1_S1752;
      end
      test_b1_S1752: begin
        IMAGE_addr <= 1736;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1753;
      end
      test_b1_S1753: begin
        IMAGE_addr <= 1737;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1724;
        test_state <= test_b1_S1754;
      end
      test_b1_S1754: begin
        IMAGE_addr <= 1738;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S1755;
      end
      test_b1_S1755: begin
        IMAGE_addr <= 1739;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 909;
        test_state <= test_b1_S1756;
      end
      test_b1_S1756: begin
        IMAGE_addr <= 1740;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 83;
        test_state <= test_b1_S1757;
      end
      test_b1_S1757: begin
        IMAGE_addr <= 1741;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 84;
        test_state <= test_b1_S1758;
      end
      test_b1_S1758: begin
        IMAGE_addr <= 1742;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 82;
        test_state <= test_b1_S1759;
      end
      test_b1_S1759: begin
        IMAGE_addr <= 1743;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 73;
        test_state <= test_b1_S1760;
      end
      test_b1_S1760: begin
        IMAGE_addr <= 1744;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 78;
        test_state <= test_b1_S1761;
      end
      test_b1_S1761: begin
        IMAGE_addr <= 1745;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 71;
        test_state <= test_b1_S1762;
      end
      test_b1_S1762: begin
        IMAGE_addr <= 1746;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 45;
        test_state <= test_b1_S1763;
      end
      test_b1_S1763: begin
        IMAGE_addr <= 1747;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 76;
        test_state <= test_b1_S1764;
      end
      test_b1_S1764: begin
        IMAGE_addr <= 1748;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 69;
        test_state <= test_b1_S1765;
      end
      test_b1_S1765: begin
        IMAGE_addr <= 1749;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 78;
        test_state <= test_b1_S1766;
      end
      test_b1_S1766: begin
        IMAGE_addr <= 1750;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 71;
        test_state <= test_b1_S1767;
      end
      test_b1_S1767: begin
        IMAGE_addr <= 1751;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 84;
        test_state <= test_b1_S1768;
      end
      test_b1_S1768: begin
        IMAGE_addr <= 1752;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 72;
        test_state <= test_b1_S1769;
      end
      test_b1_S1769: begin
        IMAGE_addr <= 1753;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1770;
      end
      test_b1_S1770: begin
        IMAGE_addr <= 1754;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1737;
        test_state <= test_b1_S1771;
      end
      test_b1_S1771: begin
        IMAGE_addr <= 1755;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S1772;
      end
      test_b1_S1772: begin
        IMAGE_addr <= 1756;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 915;
        test_state <= test_b1_S1773;
      end
      test_b1_S1773: begin
        IMAGE_addr <= 1757;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 83;
        test_state <= test_b1_S1774;
      end
      test_b1_S1774: begin
        IMAGE_addr <= 1758;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 84;
        test_state <= test_b1_S1775;
      end
      test_b1_S1775: begin
        IMAGE_addr <= 1759;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 82;
        test_state <= test_b1_S1776;
      end
      test_b1_S1776: begin
        IMAGE_addr <= 1760;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 73;
        test_state <= test_b1_S1777;
      end
      test_b1_S1777: begin
        IMAGE_addr <= 1761;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 78;
        test_state <= test_b1_S1778;
      end
      test_b1_S1778: begin
        IMAGE_addr <= 1762;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 71;
        test_state <= test_b1_S1779;
      end
      test_b1_S1779: begin
        IMAGE_addr <= 1763;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 45;
        test_state <= test_b1_S1780;
      end
      test_b1_S1780: begin
        IMAGE_addr <= 1764;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 66;
        test_state <= test_b1_S1781;
      end
      test_b1_S1781: begin
        IMAGE_addr <= 1765;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 85;
        test_state <= test_b1_S1782;
      end
      test_b1_S1782: begin
        IMAGE_addr <= 1766;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 70;
        test_state <= test_b1_S1783;
      end
      test_b1_S1783: begin
        IMAGE_addr <= 1767;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 70;
        test_state <= test_b1_S1784;
      end
      test_b1_S1784: begin
        IMAGE_addr <= 1768;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 69;
        test_state <= test_b1_S1785;
      end
      test_b1_S1785: begin
        IMAGE_addr <= 1769;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 82;
        test_state <= test_b1_S1786;
      end
      test_b1_S1786: begin
        IMAGE_addr <= 1770;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 83;
        test_state <= test_b1_S1787;
      end
      test_b1_S1787: begin
        IMAGE_addr <= 1771;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1788;
      end
      test_b1_S1788: begin
        IMAGE_addr <= 1772;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1754;
        test_state <= test_b1_S1789;
      end
      test_b1_S1789: begin
        IMAGE_addr <= 1773;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S1790;
      end
      test_b1_S1790: begin
        IMAGE_addr <= 1774;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 886;
        test_state <= test_b1_S1791;
      end
      test_b1_S1791: begin
        IMAGE_addr <= 1775;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 119;
        test_state <= test_b1_S1792;
      end
      test_b1_S1792: begin
        IMAGE_addr <= 1776;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S1793;
      end
      test_b1_S1793: begin
        IMAGE_addr <= 1777;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S1794;
      end
      test_b1_S1794: begin
        IMAGE_addr <= 1778;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 104;
        test_state <= test_b1_S1795;
      end
      test_b1_S1795: begin
        IMAGE_addr <= 1779;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 76;
        test_state <= test_b1_S1796;
      end
      test_b1_S1796: begin
        IMAGE_addr <= 1780;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S1797;
      end
      test_b1_S1797: begin
        IMAGE_addr <= 1781;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 110;
        test_state <= test_b1_S1798;
      end
      test_b1_S1798: begin
        IMAGE_addr <= 1782;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 103;
        test_state <= test_b1_S1799;
      end
      test_b1_S1799: begin
        IMAGE_addr <= 1783;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S1800;
      end
      test_b1_S1800: begin
        IMAGE_addr <= 1784;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 104;
        test_state <= test_b1_S1801;
      end
      test_b1_S1801: begin
        IMAGE_addr <= 1785;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1802;
      end
      test_b1_S1802: begin
        IMAGE_addr <= 1786;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1772;
        test_state <= test_b1_S1803;
      end
      test_b1_S1803: begin
        IMAGE_addr <= 1787;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S1804;
      end
      test_b1_S1804: begin
        IMAGE_addr <= 1788;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 286;
        test_state <= test_b1_S1805;
      end
      test_b1_S1805: begin
        IMAGE_addr <= 1789;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 119;
        test_state <= test_b1_S1806;
      end
      test_b1_S1806: begin
        IMAGE_addr <= 1790;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S1807;
      end
      test_b1_S1807: begin
        IMAGE_addr <= 1791;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S1808;
      end
      test_b1_S1808: begin
        IMAGE_addr <= 1792;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 104;
        test_state <= test_b1_S1809;
      end
      test_b1_S1809: begin
        IMAGE_addr <= 1793;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 67;
        test_state <= test_b1_S1810;
      end
      test_b1_S1810: begin
        IMAGE_addr <= 1794;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 108;
        test_state <= test_b1_S1811;
      end
      test_b1_S1811: begin
        IMAGE_addr <= 1795;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S1812;
      end
      test_b1_S1812: begin
        IMAGE_addr <= 1796;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S1813;
      end
      test_b1_S1813: begin
        IMAGE_addr <= 1797;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S1814;
      end
      test_b1_S1814: begin
        IMAGE_addr <= 1798;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1815;
      end
      test_b1_S1815: begin
        IMAGE_addr <= 1799;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1786;
        test_state <= test_b1_S1816;
      end
      test_b1_S1816: begin
        IMAGE_addr <= 1800;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S1817;
      end
      test_b1_S1817: begin
        IMAGE_addr <= 1801;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S1818;
      end
      test_b1_S1818: begin
        IMAGE_addr <= 1802;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 46;
        test_state <= test_b1_S1819;
      end
      test_b1_S1819: begin
        IMAGE_addr <= 1803;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 119;
        test_state <= test_b1_S1820;
      end
      test_b1_S1820: begin
        IMAGE_addr <= 1804;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 111;
        test_state <= test_b1_S1821;
      end
      test_b1_S1821: begin
        IMAGE_addr <= 1805;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S1822;
      end
      test_b1_S1822: begin
        IMAGE_addr <= 1806;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 100;
        test_state <= test_b1_S1823;
      end
      test_b1_S1823: begin
        IMAGE_addr <= 1807;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1824;
      end
      test_b1_S1824: begin
        IMAGE_addr <= 1808;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1799;
        test_state <= test_b1_S1825;
      end
      test_b1_S1825: begin
        IMAGE_addr <= 1809;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S1826;
      end
      test_b1_S1826: begin
        IMAGE_addr <= 1810;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 306;
        test_state <= test_b1_S1827;
      end
      test_b1_S1827: begin
        IMAGE_addr <= 1811;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 46;
        test_state <= test_b1_S1828;
      end
      test_b1_S1828: begin
        IMAGE_addr <= 1812;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 109;
        test_state <= test_b1_S1829;
      end
      test_b1_S1829: begin
        IMAGE_addr <= 1813;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S1830;
      end
      test_b1_S1830: begin
        IMAGE_addr <= 1814;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 99;
        test_state <= test_b1_S1831;
      end
      test_b1_S1831: begin
        IMAGE_addr <= 1815;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S1832;
      end
      test_b1_S1832: begin
        IMAGE_addr <= 1816;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 111;
        test_state <= test_b1_S1833;
      end
      test_b1_S1833: begin
        IMAGE_addr <= 1817;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1834;
      end
      test_b1_S1834: begin
        IMAGE_addr <= 1818;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1808;
        test_state <= test_b1_S1835;
      end
      test_b1_S1835: begin
        IMAGE_addr <= 1819;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S1836;
      end
      test_b1_S1836: begin
        IMAGE_addr <= 1820;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 310;
        test_state <= test_b1_S1837;
      end
      test_b1_S1837: begin
        IMAGE_addr <= 1821;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 46;
        test_state <= test_b1_S1838;
      end
      test_b1_S1838: begin
        IMAGE_addr <= 1822;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 100;
        test_state <= test_b1_S1839;
      end
      test_b1_S1839: begin
        IMAGE_addr <= 1823;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S1840;
      end
      test_b1_S1840: begin
        IMAGE_addr <= 1824;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S1841;
      end
      test_b1_S1841: begin
        IMAGE_addr <= 1825;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S1842;
      end
      test_b1_S1842: begin
        IMAGE_addr <= 1826;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1843;
      end
      test_b1_S1843: begin
        IMAGE_addr <= 1827;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1818;
        test_state <= test_b1_S1844;
      end
      test_b1_S1844: begin
        IMAGE_addr <= 1828;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S1845;
      end
      test_b1_S1845: begin
        IMAGE_addr <= 1829;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 323;
        test_state <= test_b1_S1846;
      end
      test_b1_S1846: begin
        IMAGE_addr <= 1830;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 46;
        test_state <= test_b1_S1847;
      end
      test_b1_S1847: begin
        IMAGE_addr <= 1831;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 112;
        test_state <= test_b1_S1848;
      end
      test_b1_S1848: begin
        IMAGE_addr <= 1832;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S1849;
      end
      test_b1_S1849: begin
        IMAGE_addr <= 1833;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S1850;
      end
      test_b1_S1850: begin
        IMAGE_addr <= 1834;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 109;
        test_state <= test_b1_S1851;
      end
      test_b1_S1851: begin
        IMAGE_addr <= 1835;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S1852;
      end
      test_b1_S1852: begin
        IMAGE_addr <= 1836;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S1853;
      end
      test_b1_S1853: begin
        IMAGE_addr <= 1837;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S1854;
      end
      test_b1_S1854: begin
        IMAGE_addr <= 1838;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 118;
        test_state <= test_b1_S1855;
      end
      test_b1_S1855: begin
        IMAGE_addr <= 1839;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S1856;
      end
      test_b1_S1856: begin
        IMAGE_addr <= 1840;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1857;
      end
      test_b1_S1857: begin
        IMAGE_addr <= 1841;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1827;
        test_state <= test_b1_S1858;
      end
      test_b1_S1858: begin
        IMAGE_addr <= 1842;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S1859;
      end
      test_b1_S1859: begin
        IMAGE_addr <= 1843;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 578;
        test_state <= test_b1_S1860;
      end
      test_b1_S1860: begin
        IMAGE_addr <= 1844;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 100;
        test_state <= test_b1_S1861;
      end
      test_b1_S1861: begin
        IMAGE_addr <= 1845;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 45;
        test_state <= test_b1_S1862;
      end
      test_b1_S1862: begin
        IMAGE_addr <= 1846;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 62;
        test_state <= test_b1_S1863;
      end
      test_b1_S1863: begin
        IMAGE_addr <= 1847;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 99;
        test_state <= test_b1_S1864;
      end
      test_b1_S1864: begin
        IMAGE_addr <= 1848;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 108;
        test_state <= test_b1_S1865;
      end
      test_b1_S1865: begin
        IMAGE_addr <= 1849;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S1866;
      end
      test_b1_S1866: begin
        IMAGE_addr <= 1850;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S1867;
      end
      test_b1_S1867: begin
        IMAGE_addr <= 1851;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S1868;
      end
      test_b1_S1868: begin
        IMAGE_addr <= 1852;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1869;
      end
      test_b1_S1869: begin
        IMAGE_addr <= 1853;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1841;
        test_state <= test_b1_S1870;
      end
      test_b1_S1870: begin
        IMAGE_addr <= 1854;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S1871;
      end
      test_b1_S1871: begin
        IMAGE_addr <= 1855;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 583;
        test_state <= test_b1_S1872;
      end
      test_b1_S1872: begin
        IMAGE_addr <= 1856;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 100;
        test_state <= test_b1_S1873;
      end
      test_b1_S1873: begin
        IMAGE_addr <= 1857;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 45;
        test_state <= test_b1_S1874;
      end
      test_b1_S1874: begin
        IMAGE_addr <= 1858;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 62;
        test_state <= test_b1_S1875;
      end
      test_b1_S1875: begin
        IMAGE_addr <= 1859;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 120;
        test_state <= test_b1_S1876;
      end
      test_b1_S1876: begin
        IMAGE_addr <= 1860;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S1877;
      end
      test_b1_S1877: begin
        IMAGE_addr <= 1861;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1878;
      end
      test_b1_S1878: begin
        IMAGE_addr <= 1862;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1853;
        test_state <= test_b1_S1879;
      end
      test_b1_S1879: begin
        IMAGE_addr <= 1863;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S1880;
      end
      test_b1_S1880: begin
        IMAGE_addr <= 1864;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 589;
        test_state <= test_b1_S1881;
      end
      test_b1_S1881: begin
        IMAGE_addr <= 1865;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 100;
        test_state <= test_b1_S1882;
      end
      test_b1_S1882: begin
        IMAGE_addr <= 1866;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 45;
        test_state <= test_b1_S1883;
      end
      test_b1_S1883: begin
        IMAGE_addr <= 1867;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 62;
        test_state <= test_b1_S1884;
      end
      test_b1_S1884: begin
        IMAGE_addr <= 1868;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 110;
        test_state <= test_b1_S1885;
      end
      test_b1_S1885: begin
        IMAGE_addr <= 1869;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S1886;
      end
      test_b1_S1886: begin
        IMAGE_addr <= 1870;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 109;
        test_state <= test_b1_S1887;
      end
      test_b1_S1887: begin
        IMAGE_addr <= 1871;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S1888;
      end
      test_b1_S1888: begin
        IMAGE_addr <= 1872;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1889;
      end
      test_b1_S1889: begin
        IMAGE_addr <= 1873;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1862;
        test_state <= test_b1_S1890;
      end
      test_b1_S1890: begin
        IMAGE_addr <= 1874;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S1891;
      end
      test_b1_S1891: begin
        IMAGE_addr <= 1875;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1110;
        test_state <= test_b1_S1892;
      end
      test_b1_S1892: begin
        IMAGE_addr <= 1876;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 98;
        test_state <= test_b1_S1893;
      end
      test_b1_S1893: begin
        IMAGE_addr <= 1877;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 111;
        test_state <= test_b1_S1894;
      end
      test_b1_S1894: begin
        IMAGE_addr <= 1878;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 111;
        test_state <= test_b1_S1895;
      end
      test_b1_S1895: begin
        IMAGE_addr <= 1879;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S1896;
      end
      test_b1_S1896: begin
        IMAGE_addr <= 1880;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1897;
      end
      test_b1_S1897: begin
        IMAGE_addr <= 1881;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1873;
        test_state <= test_b1_S1898;
      end
      test_b1_S1898: begin
        IMAGE_addr <= 1882;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S1899;
      end
      test_b1_S1899: begin
        IMAGE_addr <= 1883;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1056;
        test_state <= test_b1_S1900;
      end
      test_b1_S1900: begin
        IMAGE_addr <= 1884;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S1901;
      end
      test_b1_S1901: begin
        IMAGE_addr <= 1885;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 111;
        test_state <= test_b1_S1902;
      end
      test_b1_S1902: begin
        IMAGE_addr <= 1886;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 78;
        test_state <= test_b1_S1903;
      end
      test_b1_S1903: begin
        IMAGE_addr <= 1887;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 117;
        test_state <= test_b1_S1904;
      end
      test_b1_S1904: begin
        IMAGE_addr <= 1888;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 109;
        test_state <= test_b1_S1905;
      end
      test_b1_S1905: begin
        IMAGE_addr <= 1889;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 98;
        test_state <= test_b1_S1906;
      end
      test_b1_S1906: begin
        IMAGE_addr <= 1890;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S1907;
      end
      test_b1_S1907: begin
        IMAGE_addr <= 1891;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S1908;
      end
      test_b1_S1908: begin
        IMAGE_addr <= 1892;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1909;
      end
      test_b1_S1909: begin
        IMAGE_addr <= 1893;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1881;
        test_state <= test_b1_S1910;
      end
      test_b1_S1910: begin
        IMAGE_addr <= 1894;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S1911;
      end
      test_b1_S1911: begin
        IMAGE_addr <= 1895;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1091;
        test_state <= test_b1_S1912;
      end
      test_b1_S1912: begin
        IMAGE_addr <= 1896;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S1913;
      end
      test_b1_S1913: begin
        IMAGE_addr <= 1897;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S1914;
      end
      test_b1_S1914: begin
        IMAGE_addr <= 1898;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 78;
        test_state <= test_b1_S1915;
      end
      test_b1_S1915: begin
        IMAGE_addr <= 1899;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 117;
        test_state <= test_b1_S1916;
      end
      test_b1_S1916: begin
        IMAGE_addr <= 1900;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 109;
        test_state <= test_b1_S1917;
      end
      test_b1_S1917: begin
        IMAGE_addr <= 1901;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 98;
        test_state <= test_b1_S1918;
      end
      test_b1_S1918: begin
        IMAGE_addr <= 1902;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S1919;
      end
      test_b1_S1919: begin
        IMAGE_addr <= 1903;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S1920;
      end
      test_b1_S1920: begin
        IMAGE_addr <= 1904;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 63;
        test_state <= test_b1_S1921;
      end
      test_b1_S1921: begin
        IMAGE_addr <= 1905;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1922;
      end
      test_b1_S1922: begin
        IMAGE_addr <= 1906;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1893;
        test_state <= test_b1_S1923;
      end
      test_b1_S1923: begin
        IMAGE_addr <= 1907;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S1924;
      end
      test_b1_S1924: begin
        IMAGE_addr <= 1908;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1338;
        test_state <= test_b1_S1925;
      end
      test_b1_S1925: begin
        IMAGE_addr <= 1909;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 111;
        test_state <= test_b1_S1926;
      end
      test_b1_S1926: begin
        IMAGE_addr <= 1910;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 107;
        test_state <= test_b1_S1927;
      end
      test_b1_S1927: begin
        IMAGE_addr <= 1911;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1928;
      end
      test_b1_S1928: begin
        IMAGE_addr <= 1912;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1906;
        test_state <= test_b1_S1929;
      end
      test_b1_S1929: begin
        IMAGE_addr <= 1913;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S1930;
      end
      test_b1_S1930: begin
        IMAGE_addr <= 1914;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1385;
        test_state <= test_b1_S1931;
      end
      test_b1_S1931: begin
        IMAGE_addr <= 1915;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 108;
        test_state <= test_b1_S1932;
      end
      test_b1_S1932: begin
        IMAGE_addr <= 1916;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S1933;
      end
      test_b1_S1933: begin
        IMAGE_addr <= 1917;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S1934;
      end
      test_b1_S1934: begin
        IMAGE_addr <= 1918;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S1935;
      end
      test_b1_S1935: begin
        IMAGE_addr <= 1919;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S1936;
      end
      test_b1_S1936: begin
        IMAGE_addr <= 1920;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 110;
        test_state <= test_b1_S1937;
      end
      test_b1_S1937: begin
        IMAGE_addr <= 1921;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1938;
      end
      test_b1_S1938: begin
        IMAGE_addr <= 1922;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1912;
        test_state <= test_b1_S1939;
      end
      test_b1_S1939: begin
        IMAGE_addr <= 1923;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S1940;
      end
      test_b1_S1940: begin
        IMAGE_addr <= 1924;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 466;
        test_state <= test_b1_S1941;
      end
      test_b1_S1941: begin
        IMAGE_addr <= 1925;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 103;
        test_state <= test_b1_S1942;
      end
      test_b1_S1942: begin
        IMAGE_addr <= 1926;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S1943;
      end
      test_b1_S1943: begin
        IMAGE_addr <= 1927;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S1944;
      end
      test_b1_S1944: begin
        IMAGE_addr <= 1928;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 99;
        test_state <= test_b1_S1945;
      end
      test_b1_S1945: begin
        IMAGE_addr <= 1929;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1946;
      end
      test_b1_S1946: begin
        IMAGE_addr <= 1930;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1922;
        test_state <= test_b1_S1947;
      end
      test_b1_S1947: begin
        IMAGE_addr <= 1931;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S1948;
      end
      test_b1_S1948: begin
        IMAGE_addr <= 1932;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1232;
        test_state <= test_b1_S1949;
      end
      test_b1_S1949: begin
        IMAGE_addr <= 1933;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 102;
        test_state <= test_b1_S1950;
      end
      test_b1_S1950: begin
        IMAGE_addr <= 1934;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S1951;
      end
      test_b1_S1951: begin
        IMAGE_addr <= 1935;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 110;
        test_state <= test_b1_S1952;
      end
      test_b1_S1952: begin
        IMAGE_addr <= 1936;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 100;
        test_state <= test_b1_S1953;
      end
      test_b1_S1953: begin
        IMAGE_addr <= 1937;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1954;
      end
      test_b1_S1954: begin
        IMAGE_addr <= 1938;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1930;
        test_state <= test_b1_S1955;
      end
      test_b1_S1955: begin
        IMAGE_addr <= 1939;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S1956;
      end
      test_b1_S1956: begin
        IMAGE_addr <= 1940;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1321;
        test_state <= test_b1_S1957;
      end
      test_b1_S1957: begin
        IMAGE_addr <= 1941;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 110;
        test_state <= test_b1_S1958;
      end
      test_b1_S1958: begin
        IMAGE_addr <= 1942;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 111;
        test_state <= test_b1_S1959;
      end
      test_b1_S1959: begin
        IMAGE_addr <= 1943;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S1960;
      end
      test_b1_S1960: begin
        IMAGE_addr <= 1944;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 70;
        test_state <= test_b1_S1961;
      end
      test_b1_S1961: begin
        IMAGE_addr <= 1945;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 111;
        test_state <= test_b1_S1962;
      end
      test_b1_S1962: begin
        IMAGE_addr <= 1946;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 117;
        test_state <= test_b1_S1963;
      end
      test_b1_S1963: begin
        IMAGE_addr <= 1947;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 110;
        test_state <= test_b1_S1964;
      end
      test_b1_S1964: begin
        IMAGE_addr <= 1948;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 100;
        test_state <= test_b1_S1965;
      end
      test_b1_S1965: begin
        IMAGE_addr <= 1949;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1966;
      end
      test_b1_S1966: begin
        IMAGE_addr <= 1950;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1938;
        test_state <= test_b1_S1967;
      end
      test_b1_S1967: begin
        IMAGE_addr <= 1951;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S1968;
      end
      test_b1_S1968: begin
        IMAGE_addr <= 1952;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1310;
        test_state <= test_b1_S1969;
      end
      test_b1_S1969: begin
        IMAGE_addr <= 1953;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 60;
        test_state <= test_b1_S1970;
      end
      test_b1_S1970: begin
        IMAGE_addr <= 1954;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 110;
        test_state <= test_b1_S1971;
      end
      test_b1_S1971: begin
        IMAGE_addr <= 1955;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 111;
        test_state <= test_b1_S1972;
      end
      test_b1_S1972: begin
        IMAGE_addr <= 1956;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S1973;
      end
      test_b1_S1973: begin
        IMAGE_addr <= 1957;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 70;
        test_state <= test_b1_S1974;
      end
      test_b1_S1974: begin
        IMAGE_addr <= 1958;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 111;
        test_state <= test_b1_S1975;
      end
      test_b1_S1975: begin
        IMAGE_addr <= 1959;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 117;
        test_state <= test_b1_S1976;
      end
      test_b1_S1976: begin
        IMAGE_addr <= 1960;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 110;
        test_state <= test_b1_S1977;
      end
      test_b1_S1977: begin
        IMAGE_addr <= 1961;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 100;
        test_state <= test_b1_S1978;
      end
      test_b1_S1978: begin
        IMAGE_addr <= 1962;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 62;
        test_state <= test_b1_S1979;
      end
      test_b1_S1979: begin
        IMAGE_addr <= 1963;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1980;
      end
      test_b1_S1980: begin
        IMAGE_addr <= 1964;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1950;
        test_state <= test_b1_S1981;
      end
      test_b1_S1981: begin
        IMAGE_addr <= 1965;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S1982;
      end
      test_b1_S1982: begin
        IMAGE_addr <= 1966;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 391;
        test_state <= test_b1_S1983;
      end
      test_b1_S1983: begin
        IMAGE_addr <= 1967;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 112;
        test_state <= test_b1_S1984;
      end
      test_b1_S1984: begin
        IMAGE_addr <= 1968;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 117;
        test_state <= test_b1_S1985;
      end
      test_b1_S1985: begin
        IMAGE_addr <= 1969;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S1986;
      end
      test_b1_S1986: begin
        IMAGE_addr <= 1970;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S1987;
      end
      test_b1_S1987: begin
        IMAGE_addr <= 1971;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1988;
      end
      test_b1_S1988: begin
        IMAGE_addr <= 1972;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1964;
        test_state <= test_b1_S1989;
      end
      test_b1_S1989: begin
        IMAGE_addr <= 1973;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S1990;
      end
      test_b1_S1990: begin
        IMAGE_addr <= 1974;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 838;
        test_state <= test_b1_S1991;
      end
      test_b1_S1991: begin
        IMAGE_addr <= 1975;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 99;
        test_state <= test_b1_S1992;
      end
      test_b1_S1992: begin
        IMAGE_addr <= 1976;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 111;
        test_state <= test_b1_S1993;
      end
      test_b1_S1993: begin
        IMAGE_addr <= 1977;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 109;
        test_state <= test_b1_S1994;
      end
      test_b1_S1994: begin
        IMAGE_addr <= 1978;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 112;
        test_state <= test_b1_S1995;
      end
      test_b1_S1995: begin
        IMAGE_addr <= 1979;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S1996;
      end
      test_b1_S1996: begin
        IMAGE_addr <= 1980;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S1997;
      end
      test_b1_S1997: begin
        IMAGE_addr <= 1981;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S1998;
      end
      test_b1_S1998: begin
        IMAGE_addr <= 1982;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S1999;
      end
      test_b1_S1999: begin
        IMAGE_addr <= 1983;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1972;
        test_state <= test_b1_S2000;
      end
      test_b1_S2000: begin
        IMAGE_addr <= 1984;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S2001;
      end
      test_b1_S2001: begin
        IMAGE_addr <= 1985;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 345;
        test_state <= test_b1_S2002;
      end
      test_b1_S2002: begin
        IMAGE_addr <= 1986;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S2003;
      end
      test_b1_S2003: begin
        IMAGE_addr <= 1987;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S2004;
      end
      test_b1_S2004: begin
        IMAGE_addr <= 1988;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 100;
        test_state <= test_b1_S2005;
      end
      test_b1_S2005: begin
        IMAGE_addr <= 1989;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S2006;
      end
      test_b1_S2006: begin
        IMAGE_addr <= 1990;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S2007;
      end
      test_b1_S2007: begin
        IMAGE_addr <= 1991;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 119;
        test_state <= test_b1_S2008;
      end
      test_b1_S2008: begin
        IMAGE_addr <= 1992;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2009;
      end
      test_b1_S2009: begin
        IMAGE_addr <= 1993;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1983;
        test_state <= test_b1_S2010;
      end
      test_b1_S2010: begin
        IMAGE_addr <= 1994;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S2011;
      end
      test_b1_S2011: begin
        IMAGE_addr <= 1995;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 732;
        test_state <= test_b1_S2012;
      end
      test_b1_S2012: begin
        IMAGE_addr <= 1996;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S2013;
      end
      test_b1_S2013: begin
        IMAGE_addr <= 1997;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 102;
        test_state <= test_b1_S2014;
      end
      test_b1_S2014: begin
        IMAGE_addr <= 1998;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2015;
      end
      test_b1_S2015: begin
        IMAGE_addr <= 1999;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1993;
        test_state <= test_b1_S2016;
      end
      test_b1_S2016: begin
        IMAGE_addr <= 2000;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S2017;
      end
      test_b1_S2017: begin
        IMAGE_addr <= 2001;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 751;
        test_state <= test_b1_S2018;
      end
      test_b1_S2018: begin
        IMAGE_addr <= 2002;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S2019;
      end
      test_b1_S2019: begin
        IMAGE_addr <= 2003;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 102;
        test_state <= test_b1_S2020;
      end
      test_b1_S2020: begin
        IMAGE_addr <= 2004;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 84;
        test_state <= test_b1_S2021;
      end
      test_b1_S2021: begin
        IMAGE_addr <= 2005;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S2022;
      end
      test_b1_S2022: begin
        IMAGE_addr <= 2006;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 117;
        test_state <= test_b1_S2023;
      end
      test_b1_S2023: begin
        IMAGE_addr <= 2007;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S2024;
      end
      test_b1_S2024: begin
        IMAGE_addr <= 2008;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2025;
      end
      test_b1_S2025: begin
        IMAGE_addr <= 2009;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1999;
        test_state <= test_b1_S2026;
      end
      test_b1_S2026: begin
        IMAGE_addr <= 2010;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S2027;
      end
      test_b1_S2027: begin
        IMAGE_addr <= 2011;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 758;
        test_state <= test_b1_S2028;
      end
      test_b1_S2028: begin
        IMAGE_addr <= 2012;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S2029;
      end
      test_b1_S2029: begin
        IMAGE_addr <= 2013;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 102;
        test_state <= test_b1_S2030;
      end
      test_b1_S2030: begin
        IMAGE_addr <= 2014;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 70;
        test_state <= test_b1_S2031;
      end
      test_b1_S2031: begin
        IMAGE_addr <= 2015;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S2032;
      end
      test_b1_S2032: begin
        IMAGE_addr <= 2016;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 108;
        test_state <= test_b1_S2033;
      end
      test_b1_S2033: begin
        IMAGE_addr <= 2017;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S2034;
      end
      test_b1_S2034: begin
        IMAGE_addr <= 2018;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S2035;
      end
      test_b1_S2035: begin
        IMAGE_addr <= 2019;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2036;
      end
      test_b1_S2036: begin
        IMAGE_addr <= 2020;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2009;
        test_state <= test_b1_S2037;
      end
      test_b1_S2037: begin
        IMAGE_addr <= 2021;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S2038;
      end
      test_b1_S2038: begin
        IMAGE_addr <= 2022;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 766;
        test_state <= test_b1_S2039;
      end
      test_b1_S2039: begin
        IMAGE_addr <= 2023;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 100;
        test_state <= test_b1_S2040;
      end
      test_b1_S2040: begin
        IMAGE_addr <= 2024;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S2041;
      end
      test_b1_S2041: begin
        IMAGE_addr <= 2025;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 112;
        test_state <= test_b1_S2042;
      end
      test_b1_S2042: begin
        IMAGE_addr <= 2026;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2043;
      end
      test_b1_S2043: begin
        IMAGE_addr <= 2027;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2020;
        test_state <= test_b1_S2044;
      end
      test_b1_S2044: begin
        IMAGE_addr <= 2028;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S2045;
      end
      test_b1_S2045: begin
        IMAGE_addr <= 2029;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 774;
        test_state <= test_b1_S2046;
      end
      test_b1_S2046: begin
        IMAGE_addr <= 2030;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S2047;
      end
      test_b1_S2047: begin
        IMAGE_addr <= 2031;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S2048;
      end
      test_b1_S2048: begin
        IMAGE_addr <= 2032;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 112;
        test_state <= test_b1_S2049;
      end
      test_b1_S2049: begin
        IMAGE_addr <= 2033;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2050;
      end
      test_b1_S2050: begin
        IMAGE_addr <= 2034;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2027;
        test_state <= test_b1_S2051;
      end
      test_b1_S2051: begin
        IMAGE_addr <= 2035;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S2052;
      end
      test_b1_S2052: begin
        IMAGE_addr <= 2036;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 790;
        test_state <= test_b1_S2053;
      end
      test_b1_S2053: begin
        IMAGE_addr <= 2037;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 61;
        test_state <= test_b1_S2054;
      end
      test_b1_S2054: begin
        IMAGE_addr <= 2038;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2055;
      end
      test_b1_S2055: begin
        IMAGE_addr <= 2039;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2034;
        test_state <= test_b1_S2056;
      end
      test_b1_S2056: begin
        IMAGE_addr <= 2040;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S2057;
      end
      test_b1_S2057: begin
        IMAGE_addr <= 2041;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 798;
        test_state <= test_b1_S2058;
      end
      test_b1_S2058: begin
        IMAGE_addr <= 2042;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 60;
        test_state <= test_b1_S2059;
      end
      test_b1_S2059: begin
        IMAGE_addr <= 2043;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 62;
        test_state <= test_b1_S2060;
      end
      test_b1_S2060: begin
        IMAGE_addr <= 2044;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2061;
      end
      test_b1_S2061: begin
        IMAGE_addr <= 2045;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2039;
        test_state <= test_b1_S2062;
      end
      test_b1_S2062: begin
        IMAGE_addr <= 2046;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S2063;
      end
      test_b1_S2063: begin
        IMAGE_addr <= 2047;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 822;
        test_state <= test_b1_S2064;
      end
      test_b1_S2064: begin
        IMAGE_addr <= 2048;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 60;
        test_state <= test_b1_S2065;
      end
      test_b1_S2065: begin
        IMAGE_addr <= 2049;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2066;
      end
      test_b1_S2066: begin
        IMAGE_addr <= 2050;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2045;
        test_state <= test_b1_S2067;
      end
      test_b1_S2067: begin
        IMAGE_addr <= 2051;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S2068;
      end
      test_b1_S2068: begin
        IMAGE_addr <= 2052;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 830;
        test_state <= test_b1_S2069;
      end
      test_b1_S2069: begin
        IMAGE_addr <= 2053;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 62;
        test_state <= test_b1_S2070;
      end
      test_b1_S2070: begin
        IMAGE_addr <= 2054;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2071;
      end
      test_b1_S2071: begin
        IMAGE_addr <= 2055;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2050;
        test_state <= test_b1_S2072;
      end
      test_b1_S2072: begin
        IMAGE_addr <= 2056;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S2073;
      end
      test_b1_S2073: begin
        IMAGE_addr <= 2057;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 814;
        test_state <= test_b1_S2074;
      end
      test_b1_S2074: begin
        IMAGE_addr <= 2058;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 60;
        test_state <= test_b1_S2075;
      end
      test_b1_S2075: begin
        IMAGE_addr <= 2059;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 61;
        test_state <= test_b1_S2076;
      end
      test_b1_S2076: begin
        IMAGE_addr <= 2060;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2077;
      end
      test_b1_S2077: begin
        IMAGE_addr <= 2061;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2055;
        test_state <= test_b1_S2078;
      end
      test_b1_S2078: begin
        IMAGE_addr <= 2062;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S2079;
      end
      test_b1_S2079: begin
        IMAGE_addr <= 2063;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 806;
        test_state <= test_b1_S2080;
      end
      test_b1_S2080: begin
        IMAGE_addr <= 2064;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 62;
        test_state <= test_b1_S2081;
      end
      test_b1_S2081: begin
        IMAGE_addr <= 2065;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 61;
        test_state <= test_b1_S2082;
      end
      test_b1_S2082: begin
        IMAGE_addr <= 2066;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2083;
      end
      test_b1_S2083: begin
        IMAGE_addr <= 2067;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2061;
        test_state <= test_b1_S2084;
      end
      test_b1_S2084: begin
        IMAGE_addr <= 2068;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3283;
        test_state <= test_b1_S2085;
      end
      test_b1_S2085: begin
        IMAGE_addr <= 2069;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 229;
        test_state <= test_b1_S2086;
      end
      test_b1_S2086: begin
        IMAGE_addr <= 2070;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 59;
        test_state <= test_b1_S2087;
      end
      test_b1_S2087: begin
        IMAGE_addr <= 2071;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2088;
      end
      test_b1_S2088: begin
        IMAGE_addr <= 2072;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2067;
        test_state <= test_b1_S2089;
      end
      test_b1_S2089: begin
        IMAGE_addr <= 2073;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3283;
        test_state <= test_b1_S2090;
      end
      test_b1_S2090: begin
        IMAGE_addr <= 2074;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 222;
        test_state <= test_b1_S2091;
      end
      test_b1_S2091: begin
        IMAGE_addr <= 2075;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 59;
        test_state <= test_b1_S2092;
      end
      test_b1_S2092: begin
        IMAGE_addr <= 2076;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 59;
        test_state <= test_b1_S2093;
      end
      test_b1_S2093: begin
        IMAGE_addr <= 2077;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2094;
      end
      test_b1_S2094: begin
        IMAGE_addr <= 2078;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2072;
        test_state <= test_b1_S2095;
      end
      test_b1_S2095: begin
        IMAGE_addr <= 2079;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3283;
        test_state <= test_b1_S2096;
      end
      test_b1_S2096: begin
        IMAGE_addr <= 2080;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 273;
        test_state <= test_b1_S2097;
      end
      test_b1_S2097: begin
        IMAGE_addr <= 2081;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S2098;
      end
      test_b1_S2098: begin
        IMAGE_addr <= 2082;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S2099;
      end
      test_b1_S2099: begin
        IMAGE_addr <= 2083;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 112;
        test_state <= test_b1_S2100;
      end
      test_b1_S2100: begin
        IMAGE_addr <= 2084;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S2101;
      end
      test_b1_S2101: begin
        IMAGE_addr <= 2085;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S2102;
      end
      test_b1_S2102: begin
        IMAGE_addr <= 2086;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S2103;
      end
      test_b1_S2103: begin
        IMAGE_addr <= 2087;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2104;
      end
      test_b1_S2104: begin
        IMAGE_addr <= 2088;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2078;
        test_state <= test_b1_S2105;
      end
      test_b1_S2105: begin
        IMAGE_addr <= 2089;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3283;
        test_state <= test_b1_S2106;
      end
      test_b1_S2106: begin
        IMAGE_addr <= 2090;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 278;
        test_state <= test_b1_S2107;
      end
      test_b1_S2107: begin
        IMAGE_addr <= 2091;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S2108;
      end
      test_b1_S2108: begin
        IMAGE_addr <= 2092;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 103;
        test_state <= test_b1_S2109;
      end
      test_b1_S2109: begin
        IMAGE_addr <= 2093;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S2110;
      end
      test_b1_S2110: begin
        IMAGE_addr <= 2094;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S2111;
      end
      test_b1_S2111: begin
        IMAGE_addr <= 2095;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 110;
        test_state <= test_b1_S2112;
      end
      test_b1_S2112: begin
        IMAGE_addr <= 2096;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2113;
      end
      test_b1_S2113: begin
        IMAGE_addr <= 2097;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2088;
        test_state <= test_b1_S2114;
      end
      test_b1_S2114: begin
        IMAGE_addr <= 2098;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3283;
        test_state <= test_b1_S2115;
      end
      test_b1_S2115: begin
        IMAGE_addr <= 2099;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 266;
        test_state <= test_b1_S2116;
      end
      test_b1_S2116: begin
        IMAGE_addr <= 2100;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 48;
        test_state <= test_b1_S2117;
      end
      test_b1_S2117: begin
        IMAGE_addr <= 2101;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 59;
        test_state <= test_b1_S2118;
      end
      test_b1_S2118: begin
        IMAGE_addr <= 2102;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2119;
      end
      test_b1_S2119: begin
        IMAGE_addr <= 2103;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2097;
        test_state <= test_b1_S2120;
      end
      test_b1_S2120: begin
        IMAGE_addr <= 2104;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3283;
        test_state <= test_b1_S2121;
      end
      test_b1_S2121: begin
        IMAGE_addr <= 2105;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 252;
        test_state <= test_b1_S2122;
      end
      test_b1_S2122: begin
        IMAGE_addr <= 2106;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 112;
        test_state <= test_b1_S2123;
      end
      test_b1_S2123: begin
        IMAGE_addr <= 2107;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 117;
        test_state <= test_b1_S2124;
      end
      test_b1_S2124: begin
        IMAGE_addr <= 2108;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S2125;
      end
      test_b1_S2125: begin
        IMAGE_addr <= 2109;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 104;
        test_state <= test_b1_S2126;
      end
      test_b1_S2126: begin
        IMAGE_addr <= 2110;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2127;
      end
      test_b1_S2127: begin
        IMAGE_addr <= 2111;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2103;
        test_state <= test_b1_S2128;
      end
      test_b1_S2128: begin
        IMAGE_addr <= 2112;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3283;
        test_state <= test_b1_S2129;
      end
      test_b1_S2129: begin
        IMAGE_addr <= 2113;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 259;
        test_state <= test_b1_S2130;
      end
      test_b1_S2130: begin
        IMAGE_addr <= 2114;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 112;
        test_state <= test_b1_S2131;
      end
      test_b1_S2131: begin
        IMAGE_addr <= 2115;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 111;
        test_state <= test_b1_S2132;
      end
      test_b1_S2132: begin
        IMAGE_addr <= 2116;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 112;
        test_state <= test_b1_S2133;
      end
      test_b1_S2133: begin
        IMAGE_addr <= 2117;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2134;
      end
      test_b1_S2134: begin
        IMAGE_addr <= 2118;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2111;
        test_state <= test_b1_S2135;
      end
      test_b1_S2135: begin
        IMAGE_addr <= 2119;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 306;
        test_state <= test_b1_S2136;
      end
      test_b1_S2136: begin
        IMAGE_addr <= 2120;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 691;
        test_state <= test_b1_S2137;
      end
      test_b1_S2137: begin
        IMAGE_addr <= 2121;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 91;
        test_state <= test_b1_S2138;
      end
      test_b1_S2138: begin
        IMAGE_addr <= 2122;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2139;
      end
      test_b1_S2139: begin
        IMAGE_addr <= 2123;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2118;
        test_state <= test_b1_S2140;
      end
      test_b1_S2140: begin
        IMAGE_addr <= 2124;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 306;
        test_state <= test_b1_S2141;
      end
      test_b1_S2141: begin
        IMAGE_addr <= 2125;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 708;
        test_state <= test_b1_S2142;
      end
      test_b1_S2142: begin
        IMAGE_addr <= 2126;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 93;
        test_state <= test_b1_S2143;
      end
      test_b1_S2143: begin
        IMAGE_addr <= 2127;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2144;
      end
      test_b1_S2144: begin
        IMAGE_addr <= 2128;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2123;
        test_state <= test_b1_S2145;
      end
      test_b1_S2145: begin
        IMAGE_addr <= 2129;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 306;
        test_state <= test_b1_S2146;
      end
      test_b1_S2146: begin
        IMAGE_addr <= 2130;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 673;
        test_state <= test_b1_S2147;
      end
      test_b1_S2147: begin
        IMAGE_addr <= 2131;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 40;
        test_state <= test_b1_S2148;
      end
      test_b1_S2148: begin
        IMAGE_addr <= 2132;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2149;
      end
      test_b1_S2149: begin
        IMAGE_addr <= 2133;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2128;
        test_state <= test_b1_S2150;
      end
      test_b1_S2150: begin
        IMAGE_addr <= 2134;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 306;
        test_state <= test_b1_S2151;
      end
      test_b1_S2151: begin
        IMAGE_addr <= 2135;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 630;
        test_state <= test_b1_S2152;
      end
      test_b1_S2152: begin
        IMAGE_addr <= 2136;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 91;
        test_state <= test_b1_S2153;
      end
      test_b1_S2153: begin
        IMAGE_addr <= 2137;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 91;
        test_state <= test_b1_S2154;
      end
      test_b1_S2154: begin
        IMAGE_addr <= 2138;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2155;
      end
      test_b1_S2155: begin
        IMAGE_addr <= 2139;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2133;
        test_state <= test_b1_S2156;
      end
      test_b1_S2156: begin
        IMAGE_addr <= 2140;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 310;
        test_state <= test_b1_S2157;
      end
      test_b1_S2157: begin
        IMAGE_addr <= 2141;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S2158;
      end
      test_b1_S2158: begin
        IMAGE_addr <= 2142;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 108;
        test_state <= test_b1_S2159;
      end
      test_b1_S2159: begin
        IMAGE_addr <= 2143;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S2160;
      end
      test_b1_S2160: begin
        IMAGE_addr <= 2144;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S2161;
      end
      test_b1_S2161: begin
        IMAGE_addr <= 2145;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S2162;
      end
      test_b1_S2162: begin
        IMAGE_addr <= 2146;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2163;
      end
      test_b1_S2163: begin
        IMAGE_addr <= 2147;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2139;
        test_state <= test_b1_S2164;
      end
      test_b1_S2164: begin
        IMAGE_addr <= 2148;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 310;
        test_state <= test_b1_S2165;
      end
      test_b1_S2165: begin
        IMAGE_addr <= 2149;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S2166;
      end
      test_b1_S2166: begin
        IMAGE_addr <= 2150;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 99;
        test_state <= test_b1_S2167;
      end
      test_b1_S2167: begin
        IMAGE_addr <= 2151;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 111;
        test_state <= test_b1_S2168;
      end
      test_b1_S2168: begin
        IMAGE_addr <= 2152;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 109;
        test_state <= test_b1_S2169;
      end
      test_b1_S2169: begin
        IMAGE_addr <= 2153;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 112;
        test_state <= test_b1_S2170;
      end
      test_b1_S2170: begin
        IMAGE_addr <= 2154;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S2171;
      end
      test_b1_S2171: begin
        IMAGE_addr <= 2155;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 108;
        test_state <= test_b1_S2172;
      end
      test_b1_S2172: begin
        IMAGE_addr <= 2156;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S2173;
      end
      test_b1_S2173: begin
        IMAGE_addr <= 2157;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S2174;
      end
      test_b1_S2174: begin
        IMAGE_addr <= 2158;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2175;
      end
      test_b1_S2175: begin
        IMAGE_addr <= 2159;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2147;
        test_state <= test_b1_S2176;
      end
      test_b1_S2176: begin
        IMAGE_addr <= 2160;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 310;
        test_state <= test_b1_S2177;
      end
      test_b1_S2177: begin
        IMAGE_addr <= 2161;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1105;
        test_state <= test_b1_S2178;
      end
      test_b1_S2178: begin
        IMAGE_addr <= 2162;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 102;
        test_state <= test_b1_S2179;
      end
      test_b1_S2179: begin
        IMAGE_addr <= 2163;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 98;
        test_state <= test_b1_S2180;
      end
      test_b1_S2180: begin
        IMAGE_addr <= 2164;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2181;
      end
      test_b1_S2181: begin
        IMAGE_addr <= 2165;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2159;
        test_state <= test_b1_S2182;
      end
      test_b1_S2182: begin
        IMAGE_addr <= 2166;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 310;
        test_state <= test_b1_S2183;
      end
      test_b1_S2183: begin
        IMAGE_addr <= 2167;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1106;
        test_state <= test_b1_S2184;
      end
      test_b1_S2184: begin
        IMAGE_addr <= 2168;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 102;
        test_state <= test_b1_S2185;
      end
      test_b1_S2185: begin
        IMAGE_addr <= 2169;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 119;
        test_state <= test_b1_S2186;
      end
      test_b1_S2186: begin
        IMAGE_addr <= 2170;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2187;
      end
      test_b1_S2187: begin
        IMAGE_addr <= 2171;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2165;
        test_state <= test_b1_S2188;
      end
      test_b1_S2188: begin
        IMAGE_addr <= 2172;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 310;
        test_state <= test_b1_S2189;
      end
      test_b1_S2189: begin
        IMAGE_addr <= 2173;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1107;
        test_state <= test_b1_S2190;
      end
      test_b1_S2190: begin
        IMAGE_addr <= 2174;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 102;
        test_state <= test_b1_S2191;
      end
      test_b1_S2191: begin
        IMAGE_addr <= 2175;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 104;
        test_state <= test_b1_S2192;
      end
      test_b1_S2192: begin
        IMAGE_addr <= 2176;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2193;
      end
      test_b1_S2193: begin
        IMAGE_addr <= 2177;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2171;
        test_state <= test_b1_S2194;
      end
      test_b1_S2194: begin
        IMAGE_addr <= 2178;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 310;
        test_state <= test_b1_S2195;
      end
      test_b1_S2195: begin
        IMAGE_addr <= 2179;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1104;
        test_state <= test_b1_S2196;
      end
      test_b1_S2196: begin
        IMAGE_addr <= 2180;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 109;
        test_state <= test_b1_S2197;
      end
      test_b1_S2197: begin
        IMAGE_addr <= 2181;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S2198;
      end
      test_b1_S2198: begin
        IMAGE_addr <= 2182;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 109;
        test_state <= test_b1_S2199;
      end
      test_b1_S2199: begin
        IMAGE_addr <= 2183;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 111;
        test_state <= test_b1_S2200;
      end
      test_b1_S2200: begin
        IMAGE_addr <= 2184;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S2201;
      end
      test_b1_S2201: begin
        IMAGE_addr <= 2185;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 121;
        test_state <= test_b1_S2202;
      end
      test_b1_S2202: begin
        IMAGE_addr <= 2186;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2203;
      end
      test_b1_S2203: begin
        IMAGE_addr <= 2187;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2177;
        test_state <= test_b1_S2204;
      end
      test_b1_S2204: begin
        IMAGE_addr <= 2188;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 310;
        test_state <= test_b1_S2205;
      end
      test_b1_S2205: begin
        IMAGE_addr <= 2189;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1108;
        test_state <= test_b1_S2206;
      end
      test_b1_S2206: begin
        IMAGE_addr <= 2190;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 99;
        test_state <= test_b1_S2207;
      end
      test_b1_S2207: begin
        IMAGE_addr <= 2191;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 119;
        test_state <= test_b1_S2208;
      end
      test_b1_S2208: begin
        IMAGE_addr <= 2192;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2209;
      end
      test_b1_S2209: begin
        IMAGE_addr <= 2193;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2187;
        test_state <= test_b1_S2210;
      end
      test_b1_S2210: begin
        IMAGE_addr <= 2194;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 310;
        test_state <= test_b1_S2211;
      end
      test_b1_S2211: begin
        IMAGE_addr <= 2195;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1109;
        test_state <= test_b1_S2212;
      end
      test_b1_S2212: begin
        IMAGE_addr <= 2196;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 99;
        test_state <= test_b1_S2213;
      end
      test_b1_S2213: begin
        IMAGE_addr <= 2197;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 104;
        test_state <= test_b1_S2214;
      end
      test_b1_S2214: begin
        IMAGE_addr <= 2198;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2215;
      end
      test_b1_S2215: begin
        IMAGE_addr <= 2199;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2193;
        test_state <= test_b1_S2216;
      end
      test_b1_S2216: begin
        IMAGE_addr <= 2200;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 310;
        test_state <= test_b1_S2217;
      end
      test_b1_S2217: begin
        IMAGE_addr <= 2201;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S2218;
      end
      test_b1_S2218: begin
        IMAGE_addr <= 2202;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 104;
        test_state <= test_b1_S2219;
      end
      test_b1_S2219: begin
        IMAGE_addr <= 2203;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S2220;
      end
      test_b1_S2220: begin
        IMAGE_addr <= 2204;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S2221;
      end
      test_b1_S2221: begin
        IMAGE_addr <= 2205;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 112;
        test_state <= test_b1_S2222;
      end
      test_b1_S2222: begin
        IMAGE_addr <= 2206;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2223;
      end
      test_b1_S2223: begin
        IMAGE_addr <= 2207;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2199;
        test_state <= test_b1_S2224;
      end
      test_b1_S2224: begin
        IMAGE_addr <= 2208;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 310;
        test_state <= test_b1_S2225;
      end
      test_b1_S2225: begin
        IMAGE_addr <= 2209;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5;
        test_state <= test_b1_S2226;
      end
      test_b1_S2226: begin
        IMAGE_addr <= 2210;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 119;
        test_state <= test_b1_S2227;
      end
      test_b1_S2227: begin
        IMAGE_addr <= 2211;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 104;
        test_state <= test_b1_S2228;
      end
      test_b1_S2228: begin
        IMAGE_addr <= 2212;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S2229;
      end
      test_b1_S2229: begin
        IMAGE_addr <= 2213;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 99;
        test_state <= test_b1_S2230;
      end
      test_b1_S2230: begin
        IMAGE_addr <= 2214;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 104;
        test_state <= test_b1_S2231;
      end
      test_b1_S2231: begin
        IMAGE_addr <= 2215;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2232;
      end
      test_b1_S2232: begin
        IMAGE_addr <= 2216;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2207;
        test_state <= test_b1_S2233;
      end
      test_b1_S2233: begin
        IMAGE_addr <= 2217;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 310;
        test_state <= test_b1_S2234;
      end
      test_b1_S2234: begin
        IMAGE_addr <= 2218;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 397;
        test_state <= test_b1_S2235;
      end
      test_b1_S2235: begin
        IMAGE_addr <= 2219;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S2236;
      end
      test_b1_S2236: begin
        IMAGE_addr <= 2220;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S2237;
      end
      test_b1_S2237: begin
        IMAGE_addr <= 2221;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 109;
        test_state <= test_b1_S2238;
      end
      test_b1_S2238: begin
        IMAGE_addr <= 2222;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S2239;
      end
      test_b1_S2239: begin
        IMAGE_addr <= 2223;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 112;
        test_state <= test_b1_S2240;
      end
      test_b1_S2240: begin
        IMAGE_addr <= 2224;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 112;
        test_state <= test_b1_S2241;
      end
      test_b1_S2241: begin
        IMAGE_addr <= 2225;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S2242;
      end
      test_b1_S2242: begin
        IMAGE_addr <= 2226;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 110;
        test_state <= test_b1_S2243;
      end
      test_b1_S2243: begin
        IMAGE_addr <= 2227;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 103;
        test_state <= test_b1_S2244;
      end
      test_b1_S2244: begin
        IMAGE_addr <= 2228;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2245;
      end
      test_b1_S2245: begin
        IMAGE_addr <= 2229;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2216;
        test_state <= test_b1_S2246;
      end
      test_b1_S2246: begin
        IMAGE_addr <= 2230;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 310;
        test_state <= test_b1_S2247;
      end
      test_b1_S2247: begin
        IMAGE_addr <= 2231;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 398;
        test_state <= test_b1_S2248;
      end
      test_b1_S2248: begin
        IMAGE_addr <= 2232;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S2249;
      end
      test_b1_S2249: begin
        IMAGE_addr <= 2233;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S2250;
      end
      test_b1_S2250: begin
        IMAGE_addr <= 2234;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S2251;
      end
      test_b1_S2251: begin
        IMAGE_addr <= 2235;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 76;
        test_state <= test_b1_S2252;
      end
      test_b1_S2252: begin
        IMAGE_addr <= 2236;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S2253;
      end
      test_b1_S2253: begin
        IMAGE_addr <= 2237;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S2254;
      end
      test_b1_S2254: begin
        IMAGE_addr <= 2238;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 100;
        test_state <= test_b1_S2255;
      end
      test_b1_S2255: begin
        IMAGE_addr <= 2239;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S2256;
      end
      test_b1_S2256: begin
        IMAGE_addr <= 2240;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 110;
        test_state <= test_b1_S2257;
      end
      test_b1_S2257: begin
        IMAGE_addr <= 2241;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 103;
        test_state <= test_b1_S2258;
      end
      test_b1_S2258: begin
        IMAGE_addr <= 2242;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 63;
        test_state <= test_b1_S2259;
      end
      test_b1_S2259: begin
        IMAGE_addr <= 2243;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2260;
      end
      test_b1_S2260: begin
        IMAGE_addr <= 2244;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2229;
        test_state <= test_b1_S2261;
      end
      test_b1_S2261: begin
        IMAGE_addr <= 2245;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 310;
        test_state <= test_b1_S2262;
      end
      test_b1_S2262: begin
        IMAGE_addr <= 2246;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 925;
        test_state <= test_b1_S2263;
      end
      test_b1_S2263: begin
        IMAGE_addr <= 2247;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 98;
        test_state <= test_b1_S2264;
      end
      test_b1_S2264: begin
        IMAGE_addr <= 2248;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S2265;
      end
      test_b1_S2265: begin
        IMAGE_addr <= 2249;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S2266;
      end
      test_b1_S2266: begin
        IMAGE_addr <= 2250;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S2267;
      end
      test_b1_S2267: begin
        IMAGE_addr <= 2251;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2268;
      end
      test_b1_S2268: begin
        IMAGE_addr <= 2252;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2244;
        test_state <= test_b1_S2269;
      end
      test_b1_S2269: begin
        IMAGE_addr <= 2253;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 310;
        test_state <= test_b1_S2270;
      end
      test_b1_S2270: begin
        IMAGE_addr <= 2254;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 344;
        test_state <= test_b1_S2271;
      end
      test_b1_S2271: begin
        IMAGE_addr <= 2255;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 117;
        test_state <= test_b1_S2272;
      end
      test_b1_S2272: begin
        IMAGE_addr <= 2256;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 112;
        test_state <= test_b1_S2273;
      end
      test_b1_S2273: begin
        IMAGE_addr <= 2257;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 100;
        test_state <= test_b1_S2274;
      end
      test_b1_S2274: begin
        IMAGE_addr <= 2258;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S2275;
      end
      test_b1_S2275: begin
        IMAGE_addr <= 2259;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S2276;
      end
      test_b1_S2276: begin
        IMAGE_addr <= 2260;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S2277;
      end
      test_b1_S2277: begin
        IMAGE_addr <= 2261;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2278;
      end
      test_b1_S2278: begin
        IMAGE_addr <= 2262;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2252;
        test_state <= test_b1_S2279;
      end
      test_b1_S2279: begin
        IMAGE_addr <= 2263;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 310;
        test_state <= test_b1_S2280;
      end
      test_b1_S2280: begin
        IMAGE_addr <= 2264;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 13;
        test_state <= test_b1_S2281;
      end
      test_b1_S2281: begin
        IMAGE_addr <= 2265;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 118;
        test_state <= test_b1_S2282;
      end
      test_b1_S2282: begin
        IMAGE_addr <= 2266;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S2283;
      end
      test_b1_S2283: begin
        IMAGE_addr <= 2267;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S2284;
      end
      test_b1_S2284: begin
        IMAGE_addr <= 2268;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S2285;
      end
      test_b1_S2285: begin
        IMAGE_addr <= 2269;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S2286;
      end
      test_b1_S2286: begin
        IMAGE_addr <= 2270;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 111;
        test_state <= test_b1_S2287;
      end
      test_b1_S2287: begin
        IMAGE_addr <= 2271;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 110;
        test_state <= test_b1_S2288;
      end
      test_b1_S2288: begin
        IMAGE_addr <= 2272;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2289;
      end
      test_b1_S2289: begin
        IMAGE_addr <= 2273;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2262;
        test_state <= test_b1_S2290;
      end
      test_b1_S2290: begin
        IMAGE_addr <= 2274;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 310;
        test_state <= test_b1_S2291;
      end
      test_b1_S2291: begin
        IMAGE_addr <= 2275;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 18;
        test_state <= test_b1_S2292;
      end
      test_b1_S2292: begin
        IMAGE_addr <= 2276;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 98;
        test_state <= test_b1_S2293;
      end
      test_b1_S2293: begin
        IMAGE_addr <= 2277;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 117;
        test_state <= test_b1_S2294;
      end
      test_b1_S2294: begin
        IMAGE_addr <= 2278;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S2295;
      end
      test_b1_S2295: begin
        IMAGE_addr <= 2279;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 108;
        test_state <= test_b1_S2296;
      end
      test_b1_S2296: begin
        IMAGE_addr <= 2280;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 100;
        test_state <= test_b1_S2297;
      end
      test_b1_S2297: begin
        IMAGE_addr <= 2281;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2298;
      end
      test_b1_S2298: begin
        IMAGE_addr <= 2282;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2273;
        test_state <= test_b1_S2299;
      end
      test_b1_S2299: begin
        IMAGE_addr <= 2283;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 310;
        test_state <= test_b1_S2300;
      end
      test_b1_S2300: begin
        IMAGE_addr <= 2284;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 577;
        test_state <= test_b1_S2301;
      end
      test_b1_S2301: begin
        IMAGE_addr <= 2285;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 118;
        test_state <= test_b1_S2302;
      end
      test_b1_S2302: begin
        IMAGE_addr <= 2286;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S2303;
      end
      test_b1_S2303: begin
        IMAGE_addr <= 2287;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 99;
        test_state <= test_b1_S2304;
      end
      test_b1_S2304: begin
        IMAGE_addr <= 2288;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S2305;
      end
      test_b1_S2305: begin
        IMAGE_addr <= 2289;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 111;
        test_state <= test_b1_S2306;
      end
      test_b1_S2306: begin
        IMAGE_addr <= 2290;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S2307;
      end
      test_b1_S2307: begin
        IMAGE_addr <= 2291;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2308;
      end
      test_b1_S2308: begin
        IMAGE_addr <= 2292;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2273;
        test_state <= test_b1_S2309;
      end
      test_b1_S2309: begin
        IMAGE_addr <= 2293;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 310;
        test_state <= test_b1_S2310;
      end
      test_b1_S2310: begin
        IMAGE_addr <= 2294;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 399;
        test_state <= test_b1_S2311;
      end
      test_b1_S2311: begin
        IMAGE_addr <= 2295;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S2312;
      end
      test_b1_S2312: begin
        IMAGE_addr <= 2296;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S2313;
      end
      test_b1_S2313: begin
        IMAGE_addr <= 2297;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 98;
        test_state <= test_b1_S2314;
      end
      test_b1_S2314: begin
        IMAGE_addr <= 2298;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 65;
        test_state <= test_b1_S2315;
      end
      test_b1_S2315: begin
        IMAGE_addr <= 2299;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S2316;
      end
      test_b1_S2316: begin
        IMAGE_addr <= 2300;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 87;
        test_state <= test_b1_S2317;
      end
      test_b1_S2317: begin
        IMAGE_addr <= 2301;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 104;
        test_state <= test_b1_S2318;
      end
      test_b1_S2318: begin
        IMAGE_addr <= 2302;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S2319;
      end
      test_b1_S2319: begin
        IMAGE_addr <= 2303;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S2320;
      end
      test_b1_S2320: begin
        IMAGE_addr <= 2304;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S2321;
      end
      test_b1_S2321: begin
        IMAGE_addr <= 2305;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S2322;
      end
      test_b1_S2322: begin
        IMAGE_addr <= 2306;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 112;
        test_state <= test_b1_S2323;
      end
      test_b1_S2323: begin
        IMAGE_addr <= 2307;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S2324;
      end
      test_b1_S2324: begin
        IMAGE_addr <= 2308;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 99;
        test_state <= test_b1_S2325;
      end
      test_b1_S2325: begin
        IMAGE_addr <= 2309;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S2326;
      end
      test_b1_S2326: begin
        IMAGE_addr <= 2310;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2327;
      end
      test_b1_S2327: begin
        IMAGE_addr <= 2311;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1145;
        test_state <= test_b1_S2328;
      end
      test_b1_S2328: begin
        IMAGE_addr <= 2312;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8;
        test_state <= test_b1_S2329;
      end
      test_b1_S2329: begin
        IMAGE_addr <= 2313;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1385;
        test_state <= test_b1_S2330;
      end
      test_b1_S2330: begin
        IMAGE_addr <= 2314;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S2331;
      end
      test_b1_S2331: begin
        IMAGE_addr <= 2315;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S2332;
      end
      test_b1_S2332: begin
        IMAGE_addr <= 2316;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 118;
        test_state <= test_b1_S2333;
      end
      test_b1_S2333: begin
        IMAGE_addr <= 2317;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S2334;
      end
      test_b1_S2334: begin
        IMAGE_addr <= 2318;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2335;
      end
      test_b1_S2335: begin
        IMAGE_addr <= 2319;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 108;
        test_state <= test_b1_S2336;
      end
      test_b1_S2336: begin
        IMAGE_addr <= 2320;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2337;
      end
      test_b1_S2337: begin
        IMAGE_addr <= 2321;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 32;
        test_state <= test_b1_S2338;
      end
      test_b1_S2338: begin
        IMAGE_addr <= 2322;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S2339;
      end
      test_b1_S2339: begin
        IMAGE_addr <= 2323;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 110;
        test_state <= test_b1_S2340;
      end
      test_b1_S2340: begin
        IMAGE_addr <= 2324;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 100;
        test_state <= test_b1_S2341;
      end
      test_b1_S2341: begin
        IMAGE_addr <= 2325;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 32;
        test_state <= test_b1_S2342;
      end
      test_b1_S2342: begin
        IMAGE_addr <= 2326;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S2343;
      end
      test_b1_S2343: begin
        IMAGE_addr <= 2327;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S2344;
      end
      test_b1_S2344: begin
        IMAGE_addr <= 2328;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 118;
        test_state <= test_b1_S2345;
      end
      test_b1_S2345: begin
        IMAGE_addr <= 2329;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S2346;
      end
      test_b1_S2346: begin
        IMAGE_addr <= 2330;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 32;
        test_state <= test_b1_S2347;
      end
      test_b1_S2347: begin
        IMAGE_addr <= 2331;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 126;
        test_state <= test_b1_S2348;
      end
      test_b1_S2348: begin
        IMAGE_addr <= 2332;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 126;
        test_state <= test_b1_S2349;
      end
      test_b1_S2349: begin
        IMAGE_addr <= 2333;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 126;
        test_state <= test_b1_S2350;
      end
      test_b1_S2350: begin
        IMAGE_addr <= 2334;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 126;
        test_state <= test_b1_S2351;
      end
      test_b1_S2351: begin
        IMAGE_addr <= 2335;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 126;
        test_state <= test_b1_S2352;
      end
      test_b1_S2352: begin
        IMAGE_addr <= 2336;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 126;
        test_state <= test_b1_S2353;
      end
      test_b1_S2353: begin
        IMAGE_addr <= 2337;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 126;
        test_state <= test_b1_S2354;
      end
      test_b1_S2354: begin
        IMAGE_addr <= 2338;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 126;
        test_state <= test_b1_S2355;
      end
      test_b1_S2355: begin
        IMAGE_addr <= 2339;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 126;
        test_state <= test_b1_S2356;
      end
      test_b1_S2356: begin
        IMAGE_addr <= 2340;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 126;
        test_state <= test_b1_S2357;
      end
      test_b1_S2357: begin
        IMAGE_addr <= 2341;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 126;
        test_state <= test_b1_S2358;
      end
      test_b1_S2358: begin
        IMAGE_addr <= 2342;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 126;
        test_state <= test_b1_S2359;
      end
      test_b1_S2359: begin
        IMAGE_addr <= 2343;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 126;
        test_state <= test_b1_S2360;
      end
      test_b1_S2360: begin
        IMAGE_addr <= 2344;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 126;
        test_state <= test_b1_S2361;
      end
      test_b1_S2361: begin
        IMAGE_addr <= 2345;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 126;
        test_state <= test_b1_S2362;
      end
      test_b1_S2362: begin
        IMAGE_addr <= 2346;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 126;
        test_state <= test_b1_S2363;
      end
      test_b1_S2363: begin
        IMAGE_addr <= 2347;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 126;
        test_state <= test_b1_S2364;
      end
      test_b1_S2364: begin
        IMAGE_addr <= 2348;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 126;
        test_state <= test_b1_S2365;
      end
      test_b1_S2365: begin
        IMAGE_addr <= 2349;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 126;
        test_state <= test_b1_S2366;
      end
      test_b1_S2366: begin
        IMAGE_addr <= 2350;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 126;
        test_state <= test_b1_S2367;
      end
      test_b1_S2367: begin
        IMAGE_addr <= 2351;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 126;
        test_state <= test_b1_S2368;
      end
      test_b1_S2368: begin
        IMAGE_addr <= 2352;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 126;
        test_state <= test_b1_S2369;
      end
      test_b1_S2369: begin
        IMAGE_addr <= 2353;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 126;
        test_state <= test_b1_S2370;
      end
      test_b1_S2370: begin
        IMAGE_addr <= 2354;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 126;
        test_state <= test_b1_S2371;
      end
      test_b1_S2371: begin
        IMAGE_addr <= 2355;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 126;
        test_state <= test_b1_S2372;
      end
      test_b1_S2372: begin
        IMAGE_addr <= 2356;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 126;
        test_state <= test_b1_S2373;
      end
      test_b1_S2373: begin
        IMAGE_addr <= 2357;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 126;
        test_state <= test_b1_S2374;
      end
      test_b1_S2374: begin
        IMAGE_addr <= 2358;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 126;
        test_state <= test_b1_S2375;
      end
      test_b1_S2375: begin
        IMAGE_addr <= 2359;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 126;
        test_state <= test_b1_S2376;
      end
      test_b1_S2376: begin
        IMAGE_addr <= 2360;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 126;
        test_state <= test_b1_S2377;
      end
      test_b1_S2377: begin
        IMAGE_addr <= 2361;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 126;
        test_state <= test_b1_S2378;
      end
      test_b1_S2378: begin
        IMAGE_addr <= 2362;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 126;
        test_state <= test_b1_S2379;
      end
      test_b1_S2379: begin
        IMAGE_addr <= 2363;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 126;
        test_state <= test_b1_S2380;
      end
      test_b1_S2380: begin
        IMAGE_addr <= 2364;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 126;
        test_state <= test_b1_S2381;
      end
      test_b1_S2381: begin
        IMAGE_addr <= 2365;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 126;
        test_state <= test_b1_S2382;
      end
      test_b1_S2382: begin
        IMAGE_addr <= 2366;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 126;
        test_state <= test_b1_S2383;
      end
      test_b1_S2383: begin
        IMAGE_addr <= 2367;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 126;
        test_state <= test_b1_S2384;
      end
      test_b1_S2384: begin
        IMAGE_addr <= 2368;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 126;
        test_state <= test_b1_S2385;
      end
      test_b1_S2385: begin
        IMAGE_addr <= 2369;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 126;
        test_state <= test_b1_S2386;
      end
      test_b1_S2386: begin
        IMAGE_addr <= 2370;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 126;
        test_state <= test_b1_S2387;
      end
      test_b1_S2387: begin
        IMAGE_addr <= 2371;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 126;
        test_state <= test_b1_S2388;
      end
      test_b1_S2388: begin
        IMAGE_addr <= 2372;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 126;
        test_state <= test_b1_S2389;
      end
      test_b1_S2389: begin
        IMAGE_addr <= 2373;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 126;
        test_state <= test_b1_S2390;
      end
      test_b1_S2390: begin
        IMAGE_addr <= 2374;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 126;
        test_state <= test_b1_S2391;
      end
      test_b1_S2391: begin
        IMAGE_addr <= 2375;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 126;
        test_state <= test_b1_S2392;
      end
      test_b1_S2392: begin
        IMAGE_addr <= 2376;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 126;
        test_state <= test_b1_S2393;
      end
      test_b1_S2393: begin
        IMAGE_addr <= 2377;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 126;
        test_state <= test_b1_S2394;
      end
      test_b1_S2394: begin
        IMAGE_addr <= 2378;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 126;
        test_state <= test_b1_S2395;
      end
      test_b1_S2395: begin
        IMAGE_addr <= 2379;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 126;
        test_state <= test_b1_S2396;
      end
      test_b1_S2396: begin
        IMAGE_addr <= 2380;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 126;
        test_state <= test_b1_S2397;
      end
      test_b1_S2397: begin
        IMAGE_addr <= 2381;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 126;
        test_state <= test_b1_S2398;
      end
      test_b1_S2398: begin
        IMAGE_addr <= 2382;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 126;
        test_state <= test_b1_S2399;
      end
      test_b1_S2399: begin
        IMAGE_addr <= 2383;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 126;
        test_state <= test_b1_S2400;
      end
      test_b1_S2400: begin
        IMAGE_addr <= 2384;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 126;
        test_state <= test_b1_S2401;
      end
      test_b1_S2401: begin
        IMAGE_addr <= 2385;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 126;
        test_state <= test_b1_S2402;
      end
      test_b1_S2402: begin
        IMAGE_addr <= 2386;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 126;
        test_state <= test_b1_S2403;
      end
      test_b1_S2403: begin
        IMAGE_addr <= 2387;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 126;
        test_state <= test_b1_S2404;
      end
      test_b1_S2404: begin
        IMAGE_addr <= 2388;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 126;
        test_state <= test_b1_S2405;
      end
      test_b1_S2405: begin
        IMAGE_addr <= 2389;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 32;
        test_state <= test_b1_S2406;
      end
      test_b1_S2406: begin
        IMAGE_addr <= 2390;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2407;
      end
      test_b1_S2407: begin
        IMAGE_addr <= 2391;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2408;
      end
      test_b1_S2408: begin
        IMAGE_addr <= 2392;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2409;
      end
      test_b1_S2409: begin
        IMAGE_addr <= 2393;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2410;
      end
      test_b1_S2410: begin
        IMAGE_addr <= 2394;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2411;
      end
      test_b1_S2411: begin
        IMAGE_addr <= 2395;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2412;
      end
      test_b1_S2412: begin
        IMAGE_addr <= 2396;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2413;
      end
      test_b1_S2413: begin
        IMAGE_addr <= 2397;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2414;
      end
      test_b1_S2414: begin
        IMAGE_addr <= 2398;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2415;
      end
      test_b1_S2415: begin
        IMAGE_addr <= 2399;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2416;
      end
      test_b1_S2416: begin
        IMAGE_addr <= 2400;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2417;
      end
      test_b1_S2417: begin
        IMAGE_addr <= 2401;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2418;
      end
      test_b1_S2418: begin
        IMAGE_addr <= 2402;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2419;
      end
      test_b1_S2419: begin
        IMAGE_addr <= 2403;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2420;
      end
      test_b1_S2420: begin
        IMAGE_addr <= 2404;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2421;
      end
      test_b1_S2421: begin
        IMAGE_addr <= 2405;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2422;
      end
      test_b1_S2422: begin
        IMAGE_addr <= 2406;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2423;
      end
      test_b1_S2423: begin
        IMAGE_addr <= 2407;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2424;
      end
      test_b1_S2424: begin
        IMAGE_addr <= 2408;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2425;
      end
      test_b1_S2425: begin
        IMAGE_addr <= 2409;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2426;
      end
      test_b1_S2426: begin
        IMAGE_addr <= 2410;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2427;
      end
      test_b1_S2427: begin
        IMAGE_addr <= 2411;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2428;
      end
      test_b1_S2428: begin
        IMAGE_addr <= 2412;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2429;
      end
      test_b1_S2429: begin
        IMAGE_addr <= 2413;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2430;
      end
      test_b1_S2430: begin
        IMAGE_addr <= 2414;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2431;
      end
      test_b1_S2431: begin
        IMAGE_addr <= 2415;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2432;
      end
      test_b1_S2432: begin
        IMAGE_addr <= 2416;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2433;
      end
      test_b1_S2433: begin
        IMAGE_addr <= 2417;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2434;
      end
      test_b1_S2434: begin
        IMAGE_addr <= 2418;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2435;
      end
      test_b1_S2435: begin
        IMAGE_addr <= 2419;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2436;
      end
      test_b1_S2436: begin
        IMAGE_addr <= 2420;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2437;
      end
      test_b1_S2437: begin
        IMAGE_addr <= 2421;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2438;
      end
      test_b1_S2438: begin
        IMAGE_addr <= 2422;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2439;
      end
      test_b1_S2439: begin
        IMAGE_addr <= 2423;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2440;
      end
      test_b1_S2440: begin
        IMAGE_addr <= 2424;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2441;
      end
      test_b1_S2441: begin
        IMAGE_addr <= 2425;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2442;
      end
      test_b1_S2442: begin
        IMAGE_addr <= 2426;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2443;
      end
      test_b1_S2443: begin
        IMAGE_addr <= 2427;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2444;
      end
      test_b1_S2444: begin
        IMAGE_addr <= 2428;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2445;
      end
      test_b1_S2445: begin
        IMAGE_addr <= 2429;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2446;
      end
      test_b1_S2446: begin
        IMAGE_addr <= 2430;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2447;
      end
      test_b1_S2447: begin
        IMAGE_addr <= 2431;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2448;
      end
      test_b1_S2448: begin
        IMAGE_addr <= 2432;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2449;
      end
      test_b1_S2449: begin
        IMAGE_addr <= 2433;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2450;
      end
      test_b1_S2450: begin
        IMAGE_addr <= 2434;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2451;
      end
      test_b1_S2451: begin
        IMAGE_addr <= 2435;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2452;
      end
      test_b1_S2452: begin
        IMAGE_addr <= 2436;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2453;
      end
      test_b1_S2453: begin
        IMAGE_addr <= 2437;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2454;
      end
      test_b1_S2454: begin
        IMAGE_addr <= 2438;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2455;
      end
      test_b1_S2455: begin
        IMAGE_addr <= 2439;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2456;
      end
      test_b1_S2456: begin
        IMAGE_addr <= 2440;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2457;
      end
      test_b1_S2457: begin
        IMAGE_addr <= 2441;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2458;
      end
      test_b1_S2458: begin
        IMAGE_addr <= 2442;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2459;
      end
      test_b1_S2459: begin
        IMAGE_addr <= 2443;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2460;
      end
      test_b1_S2460: begin
        IMAGE_addr <= 2444;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2461;
      end
      test_b1_S2461: begin
        IMAGE_addr <= 2445;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2462;
      end
      test_b1_S2462: begin
        IMAGE_addr <= 2446;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2463;
      end
      test_b1_S2463: begin
        IMAGE_addr <= 2447;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2464;
      end
      test_b1_S2464: begin
        IMAGE_addr <= 2448;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2465;
      end
      test_b1_S2465: begin
        IMAGE_addr <= 2449;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2466;
      end
      test_b1_S2466: begin
        IMAGE_addr <= 2450;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2467;
      end
      test_b1_S2467: begin
        IMAGE_addr <= 2451;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2468;
      end
      test_b1_S2468: begin
        IMAGE_addr <= 2452;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2469;
      end
      test_b1_S2469: begin
        IMAGE_addr <= 2453;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2470;
      end
      test_b1_S2470: begin
        IMAGE_addr <= 2454;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2471;
      end
      test_b1_S2471: begin
        IMAGE_addr <= 2455;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2472;
      end
      test_b1_S2472: begin
        IMAGE_addr <= 2456;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2473;
      end
      test_b1_S2473: begin
        IMAGE_addr <= 2457;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2474;
      end
      test_b1_S2474: begin
        IMAGE_addr <= 2458;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2475;
      end
      test_b1_S2475: begin
        IMAGE_addr <= 2459;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2476;
      end
      test_b1_S2476: begin
        IMAGE_addr <= 2460;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2477;
      end
      test_b1_S2477: begin
        IMAGE_addr <= 2461;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2478;
      end
      test_b1_S2478: begin
        IMAGE_addr <= 2462;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2479;
      end
      test_b1_S2479: begin
        IMAGE_addr <= 2463;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2480;
      end
      test_b1_S2480: begin
        IMAGE_addr <= 2464;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2481;
      end
      test_b1_S2481: begin
        IMAGE_addr <= 2465;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2482;
      end
      test_b1_S2482: begin
        IMAGE_addr <= 2466;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2483;
      end
      test_b1_S2483: begin
        IMAGE_addr <= 2467;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2484;
      end
      test_b1_S2484: begin
        IMAGE_addr <= 2468;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2485;
      end
      test_b1_S2485: begin
        IMAGE_addr <= 2469;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2486;
      end
      test_b1_S2486: begin
        IMAGE_addr <= 2470;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2487;
      end
      test_b1_S2487: begin
        IMAGE_addr <= 2471;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2488;
      end
      test_b1_S2488: begin
        IMAGE_addr <= 2472;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2489;
      end
      test_b1_S2489: begin
        IMAGE_addr <= 2473;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2490;
      end
      test_b1_S2490: begin
        IMAGE_addr <= 2474;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2491;
      end
      test_b1_S2491: begin
        IMAGE_addr <= 2475;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2492;
      end
      test_b1_S2492: begin
        IMAGE_addr <= 2476;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2493;
      end
      test_b1_S2493: begin
        IMAGE_addr <= 2477;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2494;
      end
      test_b1_S2494: begin
        IMAGE_addr <= 2478;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2495;
      end
      test_b1_S2495: begin
        IMAGE_addr <= 2479;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2496;
      end
      test_b1_S2496: begin
        IMAGE_addr <= 2480;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2497;
      end
      test_b1_S2497: begin
        IMAGE_addr <= 2481;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2498;
      end
      test_b1_S2498: begin
        IMAGE_addr <= 2482;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2499;
      end
      test_b1_S2499: begin
        IMAGE_addr <= 2483;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2500;
      end
      test_b1_S2500: begin
        IMAGE_addr <= 2484;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2501;
      end
      test_b1_S2501: begin
        IMAGE_addr <= 2485;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2502;
      end
      test_b1_S2502: begin
        IMAGE_addr <= 2486;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2503;
      end
      test_b1_S2503: begin
        IMAGE_addr <= 2487;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2504;
      end
      test_b1_S2504: begin
        IMAGE_addr <= 2488;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2505;
      end
      test_b1_S2505: begin
        IMAGE_addr <= 2489;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2506;
      end
      test_b1_S2506: begin
        IMAGE_addr <= 2490;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2507;
      end
      test_b1_S2507: begin
        IMAGE_addr <= 2491;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2508;
      end
      test_b1_S2508: begin
        IMAGE_addr <= 2492;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2509;
      end
      test_b1_S2509: begin
        IMAGE_addr <= 2493;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2510;
      end
      test_b1_S2510: begin
        IMAGE_addr <= 2494;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2511;
      end
      test_b1_S2511: begin
        IMAGE_addr <= 2495;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2512;
      end
      test_b1_S2512: begin
        IMAGE_addr <= 2496;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2513;
      end
      test_b1_S2513: begin
        IMAGE_addr <= 2497;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2514;
      end
      test_b1_S2514: begin
        IMAGE_addr <= 2498;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2515;
      end
      test_b1_S2515: begin
        IMAGE_addr <= 2499;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2516;
      end
      test_b1_S2516: begin
        IMAGE_addr <= 2500;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2517;
      end
      test_b1_S2517: begin
        IMAGE_addr <= 2501;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2518;
      end
      test_b1_S2518: begin
        IMAGE_addr <= 2502;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2519;
      end
      test_b1_S2519: begin
        IMAGE_addr <= 2503;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2520;
      end
      test_b1_S2520: begin
        IMAGE_addr <= 2504;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2521;
      end
      test_b1_S2521: begin
        IMAGE_addr <= 2505;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2522;
      end
      test_b1_S2522: begin
        IMAGE_addr <= 2506;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2523;
      end
      test_b1_S2523: begin
        IMAGE_addr <= 2507;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2524;
      end
      test_b1_S2524: begin
        IMAGE_addr <= 2508;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2525;
      end
      test_b1_S2525: begin
        IMAGE_addr <= 2509;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2526;
      end
      test_b1_S2526: begin
        IMAGE_addr <= 2510;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2527;
      end
      test_b1_S2527: begin
        IMAGE_addr <= 2511;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2528;
      end
      test_b1_S2528: begin
        IMAGE_addr <= 2512;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2529;
      end
      test_b1_S2529: begin
        IMAGE_addr <= 2513;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2530;
      end
      test_b1_S2530: begin
        IMAGE_addr <= 2514;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2531;
      end
      test_b1_S2531: begin
        IMAGE_addr <= 2515;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2532;
      end
      test_b1_S2532: begin
        IMAGE_addr <= 2516;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2533;
      end
      test_b1_S2533: begin
        IMAGE_addr <= 2517;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2534;
      end
      test_b1_S2534: begin
        IMAGE_addr <= 2518;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2535;
      end
      test_b1_S2535: begin
        IMAGE_addr <= 2519;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2536;
      end
      test_b1_S2536: begin
        IMAGE_addr <= 2520;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2537;
      end
      test_b1_S2537: begin
        IMAGE_addr <= 2521;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2538;
      end
      test_b1_S2538: begin
        IMAGE_addr <= 2522;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2539;
      end
      test_b1_S2539: begin
        IMAGE_addr <= 2523;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2540;
      end
      test_b1_S2540: begin
        IMAGE_addr <= 2524;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2541;
      end
      test_b1_S2541: begin
        IMAGE_addr <= 2525;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2542;
      end
      test_b1_S2542: begin
        IMAGE_addr <= 2526;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2543;
      end
      test_b1_S2543: begin
        IMAGE_addr <= 2527;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2544;
      end
      test_b1_S2544: begin
        IMAGE_addr <= 2528;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2545;
      end
      test_b1_S2545: begin
        IMAGE_addr <= 2529;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2546;
      end
      test_b1_S2546: begin
        IMAGE_addr <= 2530;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2547;
      end
      test_b1_S2547: begin
        IMAGE_addr <= 2531;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2548;
      end
      test_b1_S2548: begin
        IMAGE_addr <= 2532;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2549;
      end
      test_b1_S2549: begin
        IMAGE_addr <= 2533;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2550;
      end
      test_b1_S2550: begin
        IMAGE_addr <= 2534;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2551;
      end
      test_b1_S2551: begin
        IMAGE_addr <= 2535;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2552;
      end
      test_b1_S2552: begin
        IMAGE_addr <= 2536;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2553;
      end
      test_b1_S2553: begin
        IMAGE_addr <= 2537;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2554;
      end
      test_b1_S2554: begin
        IMAGE_addr <= 2538;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2555;
      end
      test_b1_S2555: begin
        IMAGE_addr <= 2539;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2556;
      end
      test_b1_S2556: begin
        IMAGE_addr <= 2540;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2557;
      end
      test_b1_S2557: begin
        IMAGE_addr <= 2541;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2558;
      end
      test_b1_S2558: begin
        IMAGE_addr <= 2542;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2559;
      end
      test_b1_S2559: begin
        IMAGE_addr <= 2543;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2560;
      end
      test_b1_S2560: begin
        IMAGE_addr <= 2544;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2561;
      end
      test_b1_S2561: begin
        IMAGE_addr <= 2545;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2562;
      end
      test_b1_S2562: begin
        IMAGE_addr <= 2546;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2563;
      end
      test_b1_S2563: begin
        IMAGE_addr <= 2547;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2564;
      end
      test_b1_S2564: begin
        IMAGE_addr <= 2548;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2565;
      end
      test_b1_S2565: begin
        IMAGE_addr <= 2549;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2566;
      end
      test_b1_S2566: begin
        IMAGE_addr <= 2550;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2567;
      end
      test_b1_S2567: begin
        IMAGE_addr <= 2551;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2568;
      end
      test_b1_S2568: begin
        IMAGE_addr <= 2552;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2569;
      end
      test_b1_S2569: begin
        IMAGE_addr <= 2553;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2570;
      end
      test_b1_S2570: begin
        IMAGE_addr <= 2554;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2571;
      end
      test_b1_S2571: begin
        IMAGE_addr <= 2555;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2572;
      end
      test_b1_S2572: begin
        IMAGE_addr <= 2556;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2573;
      end
      test_b1_S2573: begin
        IMAGE_addr <= 2557;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2574;
      end
      test_b1_S2574: begin
        IMAGE_addr <= 2558;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2575;
      end
      test_b1_S2575: begin
        IMAGE_addr <= 2559;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2576;
      end
      test_b1_S2576: begin
        IMAGE_addr <= 2560;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2577;
      end
      test_b1_S2577: begin
        IMAGE_addr <= 2561;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2578;
      end
      test_b1_S2578: begin
        IMAGE_addr <= 2562;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2579;
      end
      test_b1_S2579: begin
        IMAGE_addr <= 2563;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2580;
      end
      test_b1_S2580: begin
        IMAGE_addr <= 2564;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2581;
      end
      test_b1_S2581: begin
        IMAGE_addr <= 2565;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2582;
      end
      test_b1_S2582: begin
        IMAGE_addr <= 2566;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2583;
      end
      test_b1_S2583: begin
        IMAGE_addr <= 2567;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2584;
      end
      test_b1_S2584: begin
        IMAGE_addr <= 2568;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2585;
      end
      test_b1_S2585: begin
        IMAGE_addr <= 2569;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2586;
      end
      test_b1_S2586: begin
        IMAGE_addr <= 2570;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2292;
        test_state <= test_b1_S2587;
      end
      test_b1_S2587: begin
        IMAGE_addr <= 2571;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S2588;
      end
      test_b1_S2588: begin
        IMAGE_addr <= 2572;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2577;
        test_state <= test_b1_S2589;
      end
      test_b1_S2589: begin
        IMAGE_addr <= 2573;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 110;
        test_state <= test_b1_S2590;
      end
      test_b1_S2590: begin
        IMAGE_addr <= 2574;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S2591;
      end
      test_b1_S2591: begin
        IMAGE_addr <= 2575;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 112;
        test_state <= test_b1_S2592;
      end
      test_b1_S2592: begin
        IMAGE_addr <= 2576;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2593;
      end
      test_b1_S2593: begin
        IMAGE_addr <= 2577;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2594;
      end
      test_b1_S2594: begin
        IMAGE_addr <= 2578;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2595;
      end
      test_b1_S2595: begin
        IMAGE_addr <= 2579;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S2596;
      end
      test_b1_S2596: begin
        IMAGE_addr <= 2580;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S2597;
      end
      test_b1_S2597: begin
        IMAGE_addr <= 2581;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S2598;
      end
      test_b1_S2598: begin
        IMAGE_addr <= 2582;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S2599;
      end
      test_b1_S2599: begin
        IMAGE_addr <= 2583;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2570;
        test_state <= test_b1_S2600;
      end
      test_b1_S2600: begin
        IMAGE_addr <= 2584;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S2601;
      end
      test_b1_S2601: begin
        IMAGE_addr <= 2585;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2590;
        test_state <= test_b1_S2602;
      end
      test_b1_S2602: begin
        IMAGE_addr <= 2586;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S2603;
      end
      test_b1_S2603: begin
        IMAGE_addr <= 2587;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 111;
        test_state <= test_b1_S2604;
      end
      test_b1_S2604: begin
        IMAGE_addr <= 2588;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S2605;
      end
      test_b1_S2605: begin
        IMAGE_addr <= 2589;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2606;
      end
      test_b1_S2606: begin
        IMAGE_addr <= 2590;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2607;
      end
      test_b1_S2607: begin
        IMAGE_addr <= 2591;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2608;
      end
      test_b1_S2608: begin
        IMAGE_addr <= 2592;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5;
        test_state <= test_b1_S2609;
      end
      test_b1_S2609: begin
        IMAGE_addr <= 2593;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S2610;
      end
      test_b1_S2610: begin
        IMAGE_addr <= 2594;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6;
        test_state <= test_b1_S2611;
      end
      test_b1_S2611: begin
        IMAGE_addr <= 2595;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S2612;
      end
      test_b1_S2612: begin
        IMAGE_addr <= 2596;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S2613;
      end
      test_b1_S2613: begin
        IMAGE_addr <= 2597;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S2614;
      end
      test_b1_S2614: begin
        IMAGE_addr <= 2598;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2583;
        test_state <= test_b1_S2615;
      end
      test_b1_S2615: begin
        IMAGE_addr <= 2599;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S2616;
      end
      test_b1_S2616: begin
        IMAGE_addr <= 2600;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2606;
        test_state <= test_b1_S2617;
      end
      test_b1_S2617: begin
        IMAGE_addr <= 2601;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S2618;
      end
      test_b1_S2618: begin
        IMAGE_addr <= 2602;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 117;
        test_state <= test_b1_S2619;
      end
      test_b1_S2619: begin
        IMAGE_addr <= 2603;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 99;
        test_state <= test_b1_S2620;
      end
      test_b1_S2620: begin
        IMAGE_addr <= 2604;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 107;
        test_state <= test_b1_S2621;
      end
      test_b1_S2621: begin
        IMAGE_addr <= 2605;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2622;
      end
      test_b1_S2622: begin
        IMAGE_addr <= 2606;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2623;
      end
      test_b1_S2623: begin
        IMAGE_addr <= 2607;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2624;
      end
      test_b1_S2624: begin
        IMAGE_addr <= 2608;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S2625;
      end
      test_b1_S2625: begin
        IMAGE_addr <= 2609;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 132;
        test_state <= test_b1_S2626;
      end
      test_b1_S2626: begin
        IMAGE_addr <= 2610;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S2627;
      end
      test_b1_S2627: begin
        IMAGE_addr <= 2611;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S2628;
      end
      test_b1_S2628: begin
        IMAGE_addr <= 2612;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2598;
        test_state <= test_b1_S2629;
      end
      test_b1_S2629: begin
        IMAGE_addr <= 2613;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S2630;
      end
      test_b1_S2630: begin
        IMAGE_addr <= 2614;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2618;
        test_state <= test_b1_S2631;
      end
      test_b1_S2631: begin
        IMAGE_addr <= 2615;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 43;
        test_state <= test_b1_S2632;
      end
      test_b1_S2632: begin
        IMAGE_addr <= 2616;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 33;
        test_state <= test_b1_S2633;
      end
      test_b1_S2633: begin
        IMAGE_addr <= 2617;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2634;
      end
      test_b1_S2634: begin
        IMAGE_addr <= 2618;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2635;
      end
      test_b1_S2635: begin
        IMAGE_addr <= 2619;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2636;
      end
      test_b1_S2636: begin
        IMAGE_addr <= 2620;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S2637;
      end
      test_b1_S2637: begin
        IMAGE_addr <= 2621;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5;
        test_state <= test_b1_S2638;
      end
      test_b1_S2638: begin
        IMAGE_addr <= 2622;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S2639;
      end
      test_b1_S2639: begin
        IMAGE_addr <= 2623;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 16;
        test_state <= test_b1_S2640;
      end
      test_b1_S2640: begin
        IMAGE_addr <= 2624;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6;
        test_state <= test_b1_S2641;
      end
      test_b1_S2641: begin
        IMAGE_addr <= 2625;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S2642;
      end
      test_b1_S2642: begin
        IMAGE_addr <= 2626;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S2643;
      end
      test_b1_S2643: begin
        IMAGE_addr <= 2627;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S2644;
      end
      test_b1_S2644: begin
        IMAGE_addr <= 2628;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2612;
        test_state <= test_b1_S2645;
      end
      test_b1_S2645: begin
        IMAGE_addr <= 2629;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S2646;
      end
      test_b1_S2646: begin
        IMAGE_addr <= 2630;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2634;
        test_state <= test_b1_S2647;
      end
      test_b1_S2647: begin
        IMAGE_addr <= 2631;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 45;
        test_state <= test_b1_S2648;
      end
      test_b1_S2648: begin
        IMAGE_addr <= 2632;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 33;
        test_state <= test_b1_S2649;
      end
      test_b1_S2649: begin
        IMAGE_addr <= 2633;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2650;
      end
      test_b1_S2650: begin
        IMAGE_addr <= 2634;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2651;
      end
      test_b1_S2651: begin
        IMAGE_addr <= 2635;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2652;
      end
      test_b1_S2652: begin
        IMAGE_addr <= 2636;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S2653;
      end
      test_b1_S2653: begin
        IMAGE_addr <= 2637;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5;
        test_state <= test_b1_S2654;
      end
      test_b1_S2654: begin
        IMAGE_addr <= 2638;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S2655;
      end
      test_b1_S2655: begin
        IMAGE_addr <= 2639;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S2656;
      end
      test_b1_S2656: begin
        IMAGE_addr <= 2640;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 17;
        test_state <= test_b1_S2657;
      end
      test_b1_S2657: begin
        IMAGE_addr <= 2641;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6;
        test_state <= test_b1_S2658;
      end
      test_b1_S2658: begin
        IMAGE_addr <= 2642;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S2659;
      end
      test_b1_S2659: begin
        IMAGE_addr <= 2643;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S2660;
      end
      test_b1_S2660: begin
        IMAGE_addr <= 2644;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S2661;
      end
      test_b1_S2661: begin
        IMAGE_addr <= 2645;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2628;
        test_state <= test_b1_S2662;
      end
      test_b1_S2662: begin
        IMAGE_addr <= 2646;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S2663;
      end
      test_b1_S2663: begin
        IMAGE_addr <= 2647;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2651;
        test_state <= test_b1_S2664;
      end
      test_b1_S2664: begin
        IMAGE_addr <= 2648;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 43;
        test_state <= test_b1_S2665;
      end
      test_b1_S2665: begin
        IMAGE_addr <= 2649;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 43;
        test_state <= test_b1_S2666;
      end
      test_b1_S2666: begin
        IMAGE_addr <= 2650;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2667;
      end
      test_b1_S2667: begin
        IMAGE_addr <= 2651;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2668;
      end
      test_b1_S2668: begin
        IMAGE_addr <= 2652;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2669;
      end
      test_b1_S2669: begin
        IMAGE_addr <= 2653;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S2670;
      end
      test_b1_S2670: begin
        IMAGE_addr <= 2654;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S2671;
      end
      test_b1_S2671: begin
        IMAGE_addr <= 2655;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S2672;
      end
      test_b1_S2672: begin
        IMAGE_addr <= 2656;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2618;
        test_state <= test_b1_S2673;
      end
      test_b1_S2673: begin
        IMAGE_addr <= 2657;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S2674;
      end
      test_b1_S2674: begin
        IMAGE_addr <= 2658;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S2675;
      end
      test_b1_S2675: begin
        IMAGE_addr <= 2659;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2645;
        test_state <= test_b1_S2676;
      end
      test_b1_S2676: begin
        IMAGE_addr <= 2660;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S2677;
      end
      test_b1_S2677: begin
        IMAGE_addr <= 2661;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2665;
        test_state <= test_b1_S2678;
      end
      test_b1_S2678: begin
        IMAGE_addr <= 2662;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 45;
        test_state <= test_b1_S2679;
      end
      test_b1_S2679: begin
        IMAGE_addr <= 2663;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 45;
        test_state <= test_b1_S2680;
      end
      test_b1_S2680: begin
        IMAGE_addr <= 2664;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2681;
      end
      test_b1_S2681: begin
        IMAGE_addr <= 2665;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2682;
      end
      test_b1_S2682: begin
        IMAGE_addr <= 2666;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2683;
      end
      test_b1_S2683: begin
        IMAGE_addr <= 2667;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S2684;
      end
      test_b1_S2684: begin
        IMAGE_addr <= 2668;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S2685;
      end
      test_b1_S2685: begin
        IMAGE_addr <= 2669;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S2686;
      end
      test_b1_S2686: begin
        IMAGE_addr <= 2670;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2634;
        test_state <= test_b1_S2687;
      end
      test_b1_S2687: begin
        IMAGE_addr <= 2671;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S2688;
      end
      test_b1_S2688: begin
        IMAGE_addr <= 2672;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S2689;
      end
      test_b1_S2689: begin
        IMAGE_addr <= 2673;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2659;
        test_state <= test_b1_S2690;
      end
      test_b1_S2690: begin
        IMAGE_addr <= 2674;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 310;
        test_state <= test_b1_S2691;
      end
      test_b1_S2691: begin
        IMAGE_addr <= 2675;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2681;
        test_state <= test_b1_S2692;
      end
      test_b1_S2692: begin
        IMAGE_addr <= 2676;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 108;
        test_state <= test_b1_S2693;
      end
      test_b1_S2693: begin
        IMAGE_addr <= 2677;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S2694;
      end
      test_b1_S2694: begin
        IMAGE_addr <= 2678;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S2695;
      end
      test_b1_S2695: begin
        IMAGE_addr <= 2679;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S2696;
      end
      test_b1_S2696: begin
        IMAGE_addr <= 2680;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2697;
      end
      test_b1_S2697: begin
        IMAGE_addr <= 2681;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8063;
        test_state <= test_b1_S2698;
      end
      test_b1_S2698: begin
        IMAGE_addr <= 2682;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8113;
        test_state <= test_b1_S2699;
      end
      test_b1_S2699: begin
        IMAGE_addr <= 2683;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2659;
        test_state <= test_b1_S2700;
      end
      test_b1_S2700: begin
        IMAGE_addr <= 2684;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S2701;
      end
      test_b1_S2701: begin
        IMAGE_addr <= 2685;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2689;
        test_state <= test_b1_S2702;
      end
      test_b1_S2702: begin
        IMAGE_addr <= 2686;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 123;
        test_state <= test_b1_S2703;
      end
      test_b1_S2703: begin
        IMAGE_addr <= 2687;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 123;
        test_state <= test_b1_S2704;
      end
      test_b1_S2704: begin
        IMAGE_addr <= 2688;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2705;
      end
      test_b1_S2705: begin
        IMAGE_addr <= 2689;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2706;
      end
      test_b1_S2706: begin
        IMAGE_addr <= 2690;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2707;
      end
      test_b1_S2707: begin
        IMAGE_addr <= 2691;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S2708;
      end
      test_b1_S2708: begin
        IMAGE_addr <= 2692;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 577;
        test_state <= test_b1_S2709;
      end
      test_b1_S2709: begin
        IMAGE_addr <= 2693;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 155;
        test_state <= test_b1_S2710;
      end
      test_b1_S2710: begin
        IMAGE_addr <= 2694;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S2711;
      end
      test_b1_S2711: begin
        IMAGE_addr <= 2695;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S2712;
      end
      test_b1_S2712: begin
        IMAGE_addr <= 2696;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S2713;
      end
      test_b1_S2713: begin
        IMAGE_addr <= 2697;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S2714;
      end
      test_b1_S2714: begin
        IMAGE_addr <= 2698;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S2715;
      end
      test_b1_S2715: begin
        IMAGE_addr <= 2699;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2681;
        test_state <= test_b1_S2716;
      end
      test_b1_S2716: begin
        IMAGE_addr <= 2700;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 197;
        test_state <= test_b1_S2717;
      end
      test_b1_S2717: begin
        IMAGE_addr <= 2701;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S2718;
      end
      test_b1_S2718: begin
        IMAGE_addr <= 2702;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S2719;
      end
      test_b1_S2719: begin
        IMAGE_addr <= 2703;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S2720;
      end
      test_b1_S2720: begin
        IMAGE_addr <= 2704;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2683;
        test_state <= test_b1_S2721;
      end
      test_b1_S2721: begin
        IMAGE_addr <= 2705;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S2722;
      end
      test_b1_S2722: begin
        IMAGE_addr <= 2706;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2720;
        test_state <= test_b1_S2723;
      end
      test_b1_S2723: begin
        IMAGE_addr <= 2707;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 45;
        test_state <= test_b1_S2724;
      end
      test_b1_S2724: begin
        IMAGE_addr <= 2708;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 45;
        test_state <= test_b1_S2725;
      end
      test_b1_S2725: begin
        IMAGE_addr <= 2709;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 45;
        test_state <= test_b1_S2726;
      end
      test_b1_S2726: begin
        IMAGE_addr <= 2710;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S2727;
      end
      test_b1_S2727: begin
        IMAGE_addr <= 2711;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S2728;
      end
      test_b1_S2728: begin
        IMAGE_addr <= 2712;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 118;
        test_state <= test_b1_S2729;
      end
      test_b1_S2729: begin
        IMAGE_addr <= 2713;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S2730;
      end
      test_b1_S2730: begin
        IMAGE_addr <= 2714;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S2731;
      end
      test_b1_S2731: begin
        IMAGE_addr <= 2715;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 108;
        test_state <= test_b1_S2732;
      end
      test_b1_S2732: begin
        IMAGE_addr <= 2716;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 45;
        test_state <= test_b1_S2733;
      end
      test_b1_S2733: begin
        IMAGE_addr <= 2717;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 45;
        test_state <= test_b1_S2734;
      end
      test_b1_S2734: begin
        IMAGE_addr <= 2718;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 45;
        test_state <= test_b1_S2735;
      end
      test_b1_S2735: begin
        IMAGE_addr <= 2719;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2736;
      end
      test_b1_S2736: begin
        IMAGE_addr <= 2720;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2737;
      end
      test_b1_S2737: begin
        IMAGE_addr <= 2721;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2738;
      end
      test_b1_S2738: begin
        IMAGE_addr <= 2722;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S2739;
      end
      test_b1_S2739: begin
        IMAGE_addr <= 2723;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 577;
        test_state <= test_b1_S2740;
      end
      test_b1_S2740: begin
        IMAGE_addr <= 2724;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 147;
        test_state <= test_b1_S2741;
      end
      test_b1_S2741: begin
        IMAGE_addr <= 2725;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S2742;
      end
      test_b1_S2742: begin
        IMAGE_addr <= 2726;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S2743;
      end
      test_b1_S2743: begin
        IMAGE_addr <= 2727;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S2744;
      end
      test_b1_S2744: begin
        IMAGE_addr <= 2728;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S2745;
      end
      test_b1_S2745: begin
        IMAGE_addr <= 2729;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2681;
        test_state <= test_b1_S2746;
      end
      test_b1_S2746: begin
        IMAGE_addr <= 2730;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 26;
        test_state <= test_b1_S2747;
      end
      test_b1_S2747: begin
        IMAGE_addr <= 2731;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S2748;
      end
      test_b1_S2748: begin
        IMAGE_addr <= 2732;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S2749;
      end
      test_b1_S2749: begin
        IMAGE_addr <= 2733;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S2750;
      end
      test_b1_S2750: begin
        IMAGE_addr <= 2734;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2704;
        test_state <= test_b1_S2751;
      end
      test_b1_S2751: begin
        IMAGE_addr <= 2735;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S2752;
      end
      test_b1_S2752: begin
        IMAGE_addr <= 2736;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2740;
        test_state <= test_b1_S2753;
      end
      test_b1_S2753: begin
        IMAGE_addr <= 2737;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 125;
        test_state <= test_b1_S2754;
      end
      test_b1_S2754: begin
        IMAGE_addr <= 2738;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 125;
        test_state <= test_b1_S2755;
      end
      test_b1_S2755: begin
        IMAGE_addr <= 2739;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2756;
      end
      test_b1_S2756: begin
        IMAGE_addr <= 2740;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2757;
      end
      test_b1_S2757: begin
        IMAGE_addr <= 2741;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2758;
      end
      test_b1_S2758: begin
        IMAGE_addr <= 2742;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S2759;
      end
      test_b1_S2759: begin
        IMAGE_addr <= 2743;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 577;
        test_state <= test_b1_S2760;
      end
      test_b1_S2760: begin
        IMAGE_addr <= 2744;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 147;
        test_state <= test_b1_S2761;
      end
      test_b1_S2761: begin
        IMAGE_addr <= 2745;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S2762;
      end
      test_b1_S2762: begin
        IMAGE_addr <= 2746;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2681;
        test_state <= test_b1_S2763;
      end
      test_b1_S2763: begin
        IMAGE_addr <= 2747;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 189;
        test_state <= test_b1_S2764;
      end
      test_b1_S2764: begin
        IMAGE_addr <= 2748;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S2765;
      end
      test_b1_S2765: begin
        IMAGE_addr <= 2749;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S2766;
      end
      test_b1_S2766: begin
        IMAGE_addr <= 2750;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 790;
        test_state <= test_b1_S2767;
      end
      test_b1_S2767: begin
        IMAGE_addr <= 2751;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S2768;
      end
      test_b1_S2768: begin
        IMAGE_addr <= 2752;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2760;
        test_state <= test_b1_S2769;
      end
      test_b1_S2769: begin
        IMAGE_addr <= 2753;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S2770;
      end
      test_b1_S2770: begin
        IMAGE_addr <= 2754;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2681;
        test_state <= test_b1_S2771;
      end
      test_b1_S2771: begin
        IMAGE_addr <= 2755;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S2772;
      end
      test_b1_S2772: begin
        IMAGE_addr <= 2756;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S2773;
      end
      test_b1_S2773: begin
        IMAGE_addr <= 2757;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S2774;
      end
      test_b1_S2774: begin
        IMAGE_addr <= 2758;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S2775;
      end
      test_b1_S2775: begin
        IMAGE_addr <= 2759;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S2776;
      end
      test_b1_S2776: begin
        IMAGE_addr <= 2760;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S2777;
      end
      test_b1_S2777: begin
        IMAGE_addr <= 2761;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2785;
        test_state <= test_b1_S2778;
      end
      test_b1_S2778: begin
        IMAGE_addr <= 2762;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S2779;
      end
      test_b1_S2779: begin
        IMAGE_addr <= 2763;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2681;
        test_state <= test_b1_S2780;
      end
      test_b1_S2780: begin
        IMAGE_addr <= 2764;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S2781;
      end
      test_b1_S2781: begin
        IMAGE_addr <= 2765;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S2782;
      end
      test_b1_S2782: begin
        IMAGE_addr <= 2766;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2782;
        test_state <= test_b1_S2783;
      end
      test_b1_S2783: begin
        IMAGE_addr <= 2767;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S2784;
      end
      test_b1_S2784: begin
        IMAGE_addr <= 2768;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S2785;
      end
      test_b1_S2785: begin
        IMAGE_addr <= 2769;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S2786;
      end
      test_b1_S2786: begin
        IMAGE_addr <= 2770;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S2787;
      end
      test_b1_S2787: begin
        IMAGE_addr <= 2771;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S2788;
      end
      test_b1_S2788: begin
        IMAGE_addr <= 2772;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S2789;
      end
      test_b1_S2789: begin
        IMAGE_addr <= 2773;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2681;
        test_state <= test_b1_S2790;
      end
      test_b1_S2790: begin
        IMAGE_addr <= 2774;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 26;
        test_state <= test_b1_S2791;
      end
      test_b1_S2791: begin
        IMAGE_addr <= 2775;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S2792;
      end
      test_b1_S2792: begin
        IMAGE_addr <= 2776;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 798;
        test_state <= test_b1_S2793;
      end
      test_b1_S2793: begin
        IMAGE_addr <= 2777;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 25;
        test_state <= test_b1_S2794;
      end
      test_b1_S2794: begin
        IMAGE_addr <= 2778;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S2795;
      end
      test_b1_S2795: begin
        IMAGE_addr <= 2779;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8;
        test_state <= test_b1_S2796;
      end
      test_b1_S2796: begin
        IMAGE_addr <= 2780;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2769;
        test_state <= test_b1_S2797;
      end
      test_b1_S2797: begin
        IMAGE_addr <= 2781;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S2798;
      end
      test_b1_S2798: begin
        IMAGE_addr <= 2782;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 183;
        test_state <= test_b1_S2799;
      end
      test_b1_S2799: begin
        IMAGE_addr <= 2783;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S2800;
      end
      test_b1_S2800: begin
        IMAGE_addr <= 2784;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S2801;
      end
      test_b1_S2801: begin
        IMAGE_addr <= 2785;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 732;
        test_state <= test_b1_S2802;
      end
      test_b1_S2802: begin
        IMAGE_addr <= 2786;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S2803;
      end
      test_b1_S2803: begin
        IMAGE_addr <= 2787;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S2804;
      end
      test_b1_S2804: begin
        IMAGE_addr <= 2788;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2734;
        test_state <= test_b1_S2805;
      end
      test_b1_S2805: begin
        IMAGE_addr <= 2789;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S2806;
      end
      test_b1_S2806: begin
        IMAGE_addr <= 2790;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2801;
        test_state <= test_b1_S2807;
      end
      test_b1_S2807: begin
        IMAGE_addr <= 2791;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 58;
        test_state <= test_b1_S2808;
      end
      test_b1_S2808: begin
        IMAGE_addr <= 2792;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 100;
        test_state <= test_b1_S2809;
      end
      test_b1_S2809: begin
        IMAGE_addr <= 2793;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S2810;
      end
      test_b1_S2810: begin
        IMAGE_addr <= 2794;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 118;
        test_state <= test_b1_S2811;
      end
      test_b1_S2811: begin
        IMAGE_addr <= 2795;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S2812;
      end
      test_b1_S2812: begin
        IMAGE_addr <= 2796;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 99;
        test_state <= test_b1_S2813;
      end
      test_b1_S2813: begin
        IMAGE_addr <= 2797;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S2814;
      end
      test_b1_S2814: begin
        IMAGE_addr <= 2798;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 111;
        test_state <= test_b1_S2815;
      end
      test_b1_S2815: begin
        IMAGE_addr <= 2799;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S2816;
      end
      test_b1_S2816: begin
        IMAGE_addr <= 2800;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2817;
      end
      test_b1_S2817: begin
        IMAGE_addr <= 2801;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2818;
      end
      test_b1_S2818: begin
        IMAGE_addr <= 2802;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2819;
      end
      test_b1_S2819: begin
        IMAGE_addr <= 2803;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S2820;
      end
      test_b1_S2820: begin
        IMAGE_addr <= 2804;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2821;
      end
      test_b1_S2821: begin
        IMAGE_addr <= 2805;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S2822;
      end
      test_b1_S2822: begin
        IMAGE_addr <= 2806;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 197;
        test_state <= test_b1_S2823;
      end
      test_b1_S2823: begin
        IMAGE_addr <= 2807;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S2824;
      end
      test_b1_S2824: begin
        IMAGE_addr <= 2808;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2825;
      end
      test_b1_S2825: begin
        IMAGE_addr <= 2809;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S2826;
      end
      test_b1_S2826: begin
        IMAGE_addr <= 2810;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S2827;
      end
      test_b1_S2827: begin
        IMAGE_addr <= 2811;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S2828;
      end
      test_b1_S2828: begin
        IMAGE_addr <= 2812;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S2829;
      end
      test_b1_S2829: begin
        IMAGE_addr <= 2813;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2788;
        test_state <= test_b1_S2830;
      end
      test_b1_S2830: begin
        IMAGE_addr <= 2814;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S2831;
      end
      test_b1_S2831: begin
        IMAGE_addr <= 2815;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2820;
        test_state <= test_b1_S2832;
      end
      test_b1_S2832: begin
        IMAGE_addr <= 2816;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 58;
        test_state <= test_b1_S2833;
      end
      test_b1_S2833: begin
        IMAGE_addr <= 2817;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S2834;
      end
      test_b1_S2834: begin
        IMAGE_addr <= 2818;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S2835;
      end
      test_b1_S2835: begin
        IMAGE_addr <= 2819;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2836;
      end
      test_b1_S2836: begin
        IMAGE_addr <= 2820;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2837;
      end
      test_b1_S2837: begin
        IMAGE_addr <= 2821;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2838;
      end
      test_b1_S2838: begin
        IMAGE_addr <= 2822;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S2839;
      end
      test_b1_S2839: begin
        IMAGE_addr <= 2823;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8;
        test_state <= test_b1_S2840;
      end
      test_b1_S2840: begin
        IMAGE_addr <= 2824;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S2841;
      end
      test_b1_S2841: begin
        IMAGE_addr <= 2825;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 197;
        test_state <= test_b1_S2842;
      end
      test_b1_S2842: begin
        IMAGE_addr <= 2826;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S2843;
      end
      test_b1_S2843: begin
        IMAGE_addr <= 2827;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S2844;
      end
      test_b1_S2844: begin
        IMAGE_addr <= 2828;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S2845;
      end
      test_b1_S2845: begin
        IMAGE_addr <= 2829;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2813;
        test_state <= test_b1_S2846;
      end
      test_b1_S2846: begin
        IMAGE_addr <= 2830;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S2847;
      end
      test_b1_S2847: begin
        IMAGE_addr <= 2831;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2841;
        test_state <= test_b1_S2848;
      end
      test_b1_S2848: begin
        IMAGE_addr <= 2832;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 100;
        test_state <= test_b1_S2849;
      end
      test_b1_S2849: begin
        IMAGE_addr <= 2833;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S2850;
      end
      test_b1_S2850: begin
        IMAGE_addr <= 2834;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 118;
        test_state <= test_b1_S2851;
      end
      test_b1_S2851: begin
        IMAGE_addr <= 2835;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S2852;
      end
      test_b1_S2852: begin
        IMAGE_addr <= 2836;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 99;
        test_state <= test_b1_S2853;
      end
      test_b1_S2853: begin
        IMAGE_addr <= 2837;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S2854;
      end
      test_b1_S2854: begin
        IMAGE_addr <= 2838;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 111;
        test_state <= test_b1_S2855;
      end
      test_b1_S2855: begin
        IMAGE_addr <= 2839;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S2856;
      end
      test_b1_S2856: begin
        IMAGE_addr <= 2840;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2857;
      end
      test_b1_S2857: begin
        IMAGE_addr <= 2841;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2858;
      end
      test_b1_S2858: begin
        IMAGE_addr <= 2842;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2859;
      end
      test_b1_S2859: begin
        IMAGE_addr <= 2843;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1239;
        test_state <= test_b1_S2860;
      end
      test_b1_S2860: begin
        IMAGE_addr <= 2844;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 25;
        test_state <= test_b1_S2861;
      end
      test_b1_S2861: begin
        IMAGE_addr <= 2845;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2801;
        test_state <= test_b1_S2862;
      end
      test_b1_S2862: begin
        IMAGE_addr <= 2846;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S2863;
      end
      test_b1_S2863: begin
        IMAGE_addr <= 2847;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S2864;
      end
      test_b1_S2864: begin
        IMAGE_addr <= 2848;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2829;
        test_state <= test_b1_S2865;
      end
      test_b1_S2865: begin
        IMAGE_addr <= 2849;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S2866;
      end
      test_b1_S2866: begin
        IMAGE_addr <= 2850;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2854;
        test_state <= test_b1_S2867;
      end
      test_b1_S2867: begin
        IMAGE_addr <= 2851;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S2868;
      end
      test_b1_S2868: begin
        IMAGE_addr <= 2852;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S2869;
      end
      test_b1_S2869: begin
        IMAGE_addr <= 2853;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2870;
      end
      test_b1_S2870: begin
        IMAGE_addr <= 2854;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2871;
      end
      test_b1_S2871: begin
        IMAGE_addr <= 2855;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2872;
      end
      test_b1_S2872: begin
        IMAGE_addr <= 2856;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1239;
        test_state <= test_b1_S2873;
      end
      test_b1_S2873: begin
        IMAGE_addr <= 2857;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 25;
        test_state <= test_b1_S2874;
      end
      test_b1_S2874: begin
        IMAGE_addr <= 2858;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2820;
        test_state <= test_b1_S2875;
      end
      test_b1_S2875: begin
        IMAGE_addr <= 2859;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S2876;
      end
      test_b1_S2876: begin
        IMAGE_addr <= 2860;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S2877;
      end
      test_b1_S2877: begin
        IMAGE_addr <= 2861;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2848;
        test_state <= test_b1_S2878;
      end
      test_b1_S2878: begin
        IMAGE_addr <= 2862;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 306;
        test_state <= test_b1_S2879;
      end
      test_b1_S2879: begin
        IMAGE_addr <= 2863;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2873;
        test_state <= test_b1_S2880;
      end
      test_b1_S2880: begin
        IMAGE_addr <= 2864;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 100;
        test_state <= test_b1_S2881;
      end
      test_b1_S2881: begin
        IMAGE_addr <= 2865;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S2882;
      end
      test_b1_S2882: begin
        IMAGE_addr <= 2866;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 102;
        test_state <= test_b1_S2883;
      end
      test_b1_S2883: begin
        IMAGE_addr <= 2867;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S2884;
      end
      test_b1_S2884: begin
        IMAGE_addr <= 2868;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 117;
        test_state <= test_b1_S2885;
      end
      test_b1_S2885: begin
        IMAGE_addr <= 2869;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 108;
        test_state <= test_b1_S2886;
      end
      test_b1_S2886: begin
        IMAGE_addr <= 2870;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S2887;
      end
      test_b1_S2887: begin
        IMAGE_addr <= 2871;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 58;
        test_state <= test_b1_S2888;
      end
      test_b1_S2888: begin
        IMAGE_addr <= 2872;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2889;
      end
      test_b1_S2889: begin
        IMAGE_addr <= 2873;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2890;
      end
      test_b1_S2890: begin
        IMAGE_addr <= 2874;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2891;
      end
      test_b1_S2891: begin
        IMAGE_addr <= 2875;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1239;
        test_state <= test_b1_S2892;
      end
      test_b1_S2892: begin
        IMAGE_addr <= 2876;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S2893;
      end
      test_b1_S2893: begin
        IMAGE_addr <= 2877;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S2894;
      end
      test_b1_S2894: begin
        IMAGE_addr <= 2878;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 16;
        test_state <= test_b1_S2895;
      end
      test_b1_S2895: begin
        IMAGE_addr <= 2879;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 213;
        test_state <= test_b1_S2896;
      end
      test_b1_S2896: begin
        IMAGE_addr <= 2880;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S2897;
      end
      test_b1_S2897: begin
        IMAGE_addr <= 2881;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S2898;
      end
      test_b1_S2898: begin
        IMAGE_addr <= 2882;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2861;
        test_state <= test_b1_S2899;
      end
      test_b1_S2899: begin
        IMAGE_addr <= 2883;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 310;
        test_state <= test_b1_S2900;
      end
      test_b1_S2900: begin
        IMAGE_addr <= 2884;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2887;
        test_state <= test_b1_S2901;
      end
      test_b1_S2901: begin
        IMAGE_addr <= 2885;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S2902;
      end
      test_b1_S2902: begin
        IMAGE_addr <= 2886;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2903;
      end
      test_b1_S2903: begin
        IMAGE_addr <= 2887;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2273;
        test_state <= test_b1_S2904;
      end
      test_b1_S2904: begin
        IMAGE_addr <= 2888;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2882;
        test_state <= test_b1_S2905;
      end
      test_b1_S2905: begin
        IMAGE_addr <= 2889;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 310;
        test_state <= test_b1_S2906;
      end
      test_b1_S2906: begin
        IMAGE_addr <= 2890;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2893;
        test_state <= test_b1_S2907;
      end
      test_b1_S2907: begin
        IMAGE_addr <= 2891;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 98;
        test_state <= test_b1_S2908;
      end
      test_b1_S2908: begin
        IMAGE_addr <= 2892;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2909;
      end
      test_b1_S2909: begin
        IMAGE_addr <= 2893;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2282;
        test_state <= test_b1_S2910;
      end
      test_b1_S2910: begin
        IMAGE_addr <= 2894;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2888;
        test_state <= test_b1_S2911;
      end
      test_b1_S2911: begin
        IMAGE_addr <= 2895;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 310;
        test_state <= test_b1_S2912;
      end
      test_b1_S2912: begin
        IMAGE_addr <= 2896;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2899;
        test_state <= test_b1_S2913;
      end
      test_b1_S2913: begin
        IMAGE_addr <= 2897;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 99;
        test_state <= test_b1_S2914;
      end
      test_b1_S2914: begin
        IMAGE_addr <= 2898;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2915;
      end
      test_b1_S2915: begin
        IMAGE_addr <= 2899;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2292;
        test_state <= test_b1_S2916;
      end
      test_b1_S2916: begin
        IMAGE_addr <= 2900;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2894;
        test_state <= test_b1_S2917;
      end
      test_b1_S2917: begin
        IMAGE_addr <= 2901;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 310;
        test_state <= test_b1_S2918;
      end
      test_b1_S2918: begin
        IMAGE_addr <= 2902;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2906;
        test_state <= test_b1_S2919;
      end
      test_b1_S2919: begin
        IMAGE_addr <= 2903;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 120;
        test_state <= test_b1_S2920;
      end
      test_b1_S2920: begin
        IMAGE_addr <= 2904;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S2921;
      end
      test_b1_S2921: begin
        IMAGE_addr <= 2905;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2922;
      end
      test_b1_S2922: begin
        IMAGE_addr <= 2906;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 577;
        test_state <= test_b1_S2923;
      end
      test_b1_S2923: begin
        IMAGE_addr <= 2907;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2900;
        test_state <= test_b1_S2924;
      end
      test_b1_S2924: begin
        IMAGE_addr <= 2908;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S2925;
      end
      test_b1_S2925: begin
        IMAGE_addr <= 2909;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2915;
        test_state <= test_b1_S2926;
      end
      test_b1_S2926: begin
        IMAGE_addr <= 2910;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S2927;
      end
      test_b1_S2927: begin
        IMAGE_addr <= 2911;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 107;
        test_state <= test_b1_S2928;
      end
      test_b1_S2928: begin
        IMAGE_addr <= 2912;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S2929;
      end
      test_b1_S2929: begin
        IMAGE_addr <= 2913;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 109;
        test_state <= test_b1_S2930;
      end
      test_b1_S2930: begin
        IMAGE_addr <= 2914;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2931;
      end
      test_b1_S2931: begin
        IMAGE_addr <= 2915;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S2932;
      end
      test_b1_S2932: begin
        IMAGE_addr <= 2916;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S2933;
      end
      test_b1_S2933: begin
        IMAGE_addr <= 2917;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S2934;
      end
      test_b1_S2934: begin
        IMAGE_addr <= 2918;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 132;
        test_state <= test_b1_S2935;
      end
      test_b1_S2935: begin
        IMAGE_addr <= 2919;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 132;
        test_state <= test_b1_S2936;
      end
      test_b1_S2936: begin
        IMAGE_addr <= 2920;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 583;
        test_state <= test_b1_S2937;
      end
      test_b1_S2937: begin
        IMAGE_addr <= 2921;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S2938;
      end
      test_b1_S2938: begin
        IMAGE_addr <= 2922;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 790;
        test_state <= test_b1_S2939;
      end
      test_b1_S2939: begin
        IMAGE_addr <= 2923;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S2940;
      end
      test_b1_S2940: begin
        IMAGE_addr <= 2924;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2929;
        test_state <= test_b1_S2941;
      end
      test_b1_S2941: begin
        IMAGE_addr <= 2925;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2577;
        test_state <= test_b1_S2942;
      end
      test_b1_S2942: begin
        IMAGE_addr <= 2926;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S2943;
      end
      test_b1_S2943: begin
        IMAGE_addr <= 2927;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2944;
      end
      test_b1_S2944: begin
        IMAGE_addr <= 2928;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S2945;
      end
      test_b1_S2945: begin
        IMAGE_addr <= 2929;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 751;
        test_state <= test_b1_S2946;
      end
      test_b1_S2946: begin
        IMAGE_addr <= 2930;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 25;
        test_state <= test_b1_S2947;
      end
      test_b1_S2947: begin
        IMAGE_addr <= 2931;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8;
        test_state <= test_b1_S2948;
      end
      test_b1_S2948: begin
        IMAGE_addr <= 2932;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2917;
        test_state <= test_b1_S2949;
      end
      test_b1_S2949: begin
        IMAGE_addr <= 2933;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S2950;
      end
      test_b1_S2950: begin
        IMAGE_addr <= 2934;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S2951;
      end
      test_b1_S2951: begin
        IMAGE_addr <= 2935;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2907;
        test_state <= test_b1_S2952;
      end
      test_b1_S2952: begin
        IMAGE_addr <= 2936;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S2953;
      end
      test_b1_S2953: begin
        IMAGE_addr <= 2937;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2949;
        test_state <= test_b1_S2954;
      end
      test_b1_S2954: begin
        IMAGE_addr <= 2938;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 103;
        test_state <= test_b1_S2955;
      end
      test_b1_S2955: begin
        IMAGE_addr <= 2939;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S2956;
      end
      test_b1_S2956: begin
        IMAGE_addr <= 2940;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S2957;
      end
      test_b1_S2957: begin
        IMAGE_addr <= 2941;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 72;
        test_state <= test_b1_S2958;
      end
      test_b1_S2958: begin
        IMAGE_addr <= 2942;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S2959;
      end
      test_b1_S2959: begin
        IMAGE_addr <= 2943;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S2960;
      end
      test_b1_S2960: begin
        IMAGE_addr <= 2944;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 100;
        test_state <= test_b1_S2961;
      end
      test_b1_S2961: begin
        IMAGE_addr <= 2945;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S2962;
      end
      test_b1_S2962: begin
        IMAGE_addr <= 2946;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S2963;
      end
      test_b1_S2963: begin
        IMAGE_addr <= 2947;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S2964;
      end
      test_b1_S2964: begin
        IMAGE_addr <= 2948;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2965;
      end
      test_b1_S2965: begin
        IMAGE_addr <= 2949;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S2966;
      end
      test_b1_S2966: begin
        IMAGE_addr <= 2950;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2906;
        test_state <= test_b1_S2967;
      end
      test_b1_S2967: begin
        IMAGE_addr <= 2951;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S2968;
      end
      test_b1_S2968: begin
        IMAGE_addr <= 2952;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S2969;
      end
      test_b1_S2969: begin
        IMAGE_addr <= 2953;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2970;
      end
      test_b1_S2970: begin
        IMAGE_addr <= 2954;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S2971;
      end
      test_b1_S2971: begin
        IMAGE_addr <= 2955;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2887;
        test_state <= test_b1_S2972;
      end
      test_b1_S2972: begin
        IMAGE_addr <= 2956;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S2973;
      end
      test_b1_S2973: begin
        IMAGE_addr <= 2957;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S2974;
      end
      test_b1_S2974: begin
        IMAGE_addr <= 2958;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2975;
      end
      test_b1_S2975: begin
        IMAGE_addr <= 2959;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S2976;
      end
      test_b1_S2976: begin
        IMAGE_addr <= 2960;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2893;
        test_state <= test_b1_S2977;
      end
      test_b1_S2977: begin
        IMAGE_addr <= 2961;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S2978;
      end
      test_b1_S2978: begin
        IMAGE_addr <= 2962;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S2979;
      end
      test_b1_S2979: begin
        IMAGE_addr <= 2963;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S2980;
      end
      test_b1_S2980: begin
        IMAGE_addr <= 2964;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S2981;
      end
      test_b1_S2981: begin
        IMAGE_addr <= 2965;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2899;
        test_state <= test_b1_S2982;
      end
      test_b1_S2982: begin
        IMAGE_addr <= 2966;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S2983;
      end
      test_b1_S2983: begin
        IMAGE_addr <= 2967;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S2984;
      end
      test_b1_S2984: begin
        IMAGE_addr <= 2968;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S2985;
      end
      test_b1_S2985: begin
        IMAGE_addr <= 2969;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S2986;
      end
      test_b1_S2986: begin
        IMAGE_addr <= 2970;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 25;
        test_state <= test_b1_S2987;
      end
      test_b1_S2987: begin
        IMAGE_addr <= 2971;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S2988;
      end
      test_b1_S2988: begin
        IMAGE_addr <= 2972;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 583;
        test_state <= test_b1_S2989;
      end
      test_b1_S2989: begin
        IMAGE_addr <= 2973;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S2990;
      end
      test_b1_S2990: begin
        IMAGE_addr <= 2974;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S2991;
      end
      test_b1_S2991: begin
        IMAGE_addr <= 2975;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2906;
        test_state <= test_b1_S2992;
      end
      test_b1_S2992: begin
        IMAGE_addr <= 2976;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S2993;
      end
      test_b1_S2993: begin
        IMAGE_addr <= 2977;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 790;
        test_state <= test_b1_S2994;
      end
      test_b1_S2994: begin
        IMAGE_addr <= 2978;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S2995;
      end
      test_b1_S2995: begin
        IMAGE_addr <= 2979;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2991;
        test_state <= test_b1_S2996;
      end
      test_b1_S2996: begin
        IMAGE_addr <= 2980;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S2997;
      end
      test_b1_S2997: begin
        IMAGE_addr <= 2981;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S2998;
      end
      test_b1_S2998: begin
        IMAGE_addr <= 2982;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2893;
        test_state <= test_b1_S2999;
      end
      test_b1_S2999: begin
        IMAGE_addr <= 2983;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S3000;
      end
      test_b1_S3000: begin
        IMAGE_addr <= 2984;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S3001;
      end
      test_b1_S3001: begin
        IMAGE_addr <= 2985;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S3002;
      end
      test_b1_S3002: begin
        IMAGE_addr <= 2986;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2887;
        test_state <= test_b1_S3003;
      end
      test_b1_S3003: begin
        IMAGE_addr <= 2987;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S3004;
      end
      test_b1_S3004: begin
        IMAGE_addr <= 2988;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S3005;
      end
      test_b1_S3005: begin
        IMAGE_addr <= 2989;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3006;
      end
      test_b1_S3006: begin
        IMAGE_addr <= 2990;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3007;
      end
      test_b1_S3007: begin
        IMAGE_addr <= 2991;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S3008;
      end
      test_b1_S3008: begin
        IMAGE_addr <= 2992;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2996;
        test_state <= test_b1_S3009;
      end
      test_b1_S3009: begin
        IMAGE_addr <= 2993;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S3010;
      end
      test_b1_S3010: begin
        IMAGE_addr <= 2994;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4294967295;
        test_state <= test_b1_S3011;
      end
      test_b1_S3011: begin
        IMAGE_addr <= 2995;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3012;
      end
      test_b1_S3012: begin
        IMAGE_addr <= 2996;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 732;
        test_state <= test_b1_S3013;
      end
      test_b1_S3013: begin
        IMAGE_addr <= 2997;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 25;
        test_state <= test_b1_S3014;
      end
      test_b1_S3014: begin
        IMAGE_addr <= 2998;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S3015;
      end
      test_b1_S3015: begin
        IMAGE_addr <= 2999;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S3016;
      end
      test_b1_S3016: begin
        IMAGE_addr <= 3000;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S3017;
      end
      test_b1_S3017: begin
        IMAGE_addr <= 3001;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2899;
        test_state <= test_b1_S3018;
      end
      test_b1_S3018: begin
        IMAGE_addr <= 3002;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S3019;
      end
      test_b1_S3019: begin
        IMAGE_addr <= 3003;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8;
        test_state <= test_b1_S3020;
      end
      test_b1_S3020: begin
        IMAGE_addr <= 3004;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2969;
        test_state <= test_b1_S3021;
      end
      test_b1_S3021: begin
        IMAGE_addr <= 3005;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3022;
      end
      test_b1_S3022: begin
        IMAGE_addr <= 3006;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3023;
      end
      test_b1_S3023: begin
        IMAGE_addr <= 3007;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2935;
        test_state <= test_b1_S3024;
      end
      test_b1_S3024: begin
        IMAGE_addr <= 3008;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S3025;
      end
      test_b1_S3025: begin
        IMAGE_addr <= 3009;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3017;
        test_state <= test_b1_S3026;
      end
      test_b1_S3026: begin
        IMAGE_addr <= 3010;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 60;
        test_state <= test_b1_S3027;
      end
      test_b1_S3027: begin
        IMAGE_addr <= 3011;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 104;
        test_state <= test_b1_S3028;
      end
      test_b1_S3028: begin
        IMAGE_addr <= 3012;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S3029;
      end
      test_b1_S3029: begin
        IMAGE_addr <= 3013;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 100;
        test_state <= test_b1_S3030;
      end
      test_b1_S3030: begin
        IMAGE_addr <= 3014;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S3031;
      end
      test_b1_S3031: begin
        IMAGE_addr <= 3015;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 62;
        test_state <= test_b1_S3032;
      end
      test_b1_S3032: begin
        IMAGE_addr <= 3016;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3033;
      end
      test_b1_S3033: begin
        IMAGE_addr <= 3017;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2949;
        test_state <= test_b1_S3034;
      end
      test_b1_S3034: begin
        IMAGE_addr <= 3018;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S3035;
      end
      test_b1_S3035: begin
        IMAGE_addr <= 3019;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2893;
        test_state <= test_b1_S3036;
      end
      test_b1_S3036: begin
        IMAGE_addr <= 3020;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S3037;
      end
      test_b1_S3037: begin
        IMAGE_addr <= 3021;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 25;
        test_state <= test_b1_S3038;
      end
      test_b1_S3038: begin
        IMAGE_addr <= 3022;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S3039;
      end
      test_b1_S3039: begin
        IMAGE_addr <= 3023;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S3040;
      end
      test_b1_S3040: begin
        IMAGE_addr <= 3024;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2887;
        test_state <= test_b1_S3041;
      end
      test_b1_S3041: begin
        IMAGE_addr <= 3025;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S3042;
      end
      test_b1_S3042: begin
        IMAGE_addr <= 3026;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S3043;
      end
      test_b1_S3043: begin
        IMAGE_addr <= 3027;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2899;
        test_state <= test_b1_S3044;
      end
      test_b1_S3044: begin
        IMAGE_addr <= 3028;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S3045;
      end
      test_b1_S3045: begin
        IMAGE_addr <= 3029;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S3046;
      end
      test_b1_S3046: begin
        IMAGE_addr <= 3030;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3047;
      end
      test_b1_S3047: begin
        IMAGE_addr <= 3031;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3048;
      end
      test_b1_S3048: begin
        IMAGE_addr <= 3032;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2861;
        test_state <= test_b1_S3049;
      end
      test_b1_S3049: begin
        IMAGE_addr <= 3033;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S3050;
      end
      test_b1_S3050: begin
        IMAGE_addr <= 3034;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3038;
        test_state <= test_b1_S3051;
      end
      test_b1_S3051: begin
        IMAGE_addr <= 3035;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 100;
        test_state <= test_b1_S3052;
      end
      test_b1_S3052: begin
        IMAGE_addr <= 3036;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 39;
        test_state <= test_b1_S3053;
      end
      test_b1_S3053: begin
        IMAGE_addr <= 3037;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3054;
      end
      test_b1_S3054: begin
        IMAGE_addr <= 3038;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3055;
      end
      test_b1_S3055: begin
        IMAGE_addr <= 3039;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3056;
      end
      test_b1_S3056: begin
        IMAGE_addr <= 3040;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1239;
        test_state <= test_b1_S3057;
      end
      test_b1_S3057: begin
        IMAGE_addr <= 3041;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S3058;
      end
      test_b1_S3058: begin
        IMAGE_addr <= 3042;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S3059;
      end
      test_b1_S3059: begin
        IMAGE_addr <= 3043;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5;
        test_state <= test_b1_S3060;
      end
      test_b1_S3060: begin
        IMAGE_addr <= 3044;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S3061;
      end
      test_b1_S3061: begin
        IMAGE_addr <= 3045;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3062;
      end
      test_b1_S3062: begin
        IMAGE_addr <= 3046;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3063;
      end
      test_b1_S3063: begin
        IMAGE_addr <= 3047;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3032;
        test_state <= test_b1_S3064;
      end
      test_b1_S3064: begin
        IMAGE_addr <= 3048;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S3065;
      end
      test_b1_S3065: begin
        IMAGE_addr <= 3049;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3056;
        test_state <= test_b1_S3066;
      end
      test_b1_S3066: begin
        IMAGE_addr <= 3050;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 120;
        test_state <= test_b1_S3067;
      end
      test_b1_S3067: begin
        IMAGE_addr <= 3051;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S3068;
      end
      test_b1_S3068: begin
        IMAGE_addr <= 3052;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 45;
        test_state <= test_b1_S3069;
      end
      test_b1_S3069: begin
        IMAGE_addr <= 3053;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 62;
        test_state <= test_b1_S3070;
      end
      test_b1_S3070: begin
        IMAGE_addr <= 3054;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 100;
        test_state <= test_b1_S3071;
      end
      test_b1_S3071: begin
        IMAGE_addr <= 3055;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3072;
      end
      test_b1_S3072: begin
        IMAGE_addr <= 3056;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8;
        test_state <= test_b1_S3073;
      end
      test_b1_S3073: begin
        IMAGE_addr <= 3057;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5522;
        test_state <= test_b1_S3074;
      end
      test_b1_S3074: begin
        IMAGE_addr <= 3058;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S3075;
      end
      test_b1_S3075: begin
        IMAGE_addr <= 3059;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2915;
        test_state <= test_b1_S3076;
      end
      test_b1_S3076: begin
        IMAGE_addr <= 3060;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 132;
        test_state <= test_b1_S3077;
      end
      test_b1_S3077: begin
        IMAGE_addr <= 3061;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 132;
        test_state <= test_b1_S3078;
      end
      test_b1_S3078: begin
        IMAGE_addr <= 3062;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 790;
        test_state <= test_b1_S3079;
      end
      test_b1_S3079: begin
        IMAGE_addr <= 3063;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S3080;
      end
      test_b1_S3080: begin
        IMAGE_addr <= 3064;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3067;
        test_state <= test_b1_S3081;
      end
      test_b1_S3081: begin
        IMAGE_addr <= 3065;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 17;
        test_state <= test_b1_S3082;
      end
      test_b1_S3082: begin
        IMAGE_addr <= 3066;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3083;
      end
      test_b1_S3083: begin
        IMAGE_addr <= 3067;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S3084;
      end
      test_b1_S3084: begin
        IMAGE_addr <= 3068;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3071;
        test_state <= test_b1_S3085;
      end
      test_b1_S3085: begin
        IMAGE_addr <= 3069;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2577;
        test_state <= test_b1_S3086;
      end
      test_b1_S3086: begin
        IMAGE_addr <= 3070;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3087;
      end
      test_b1_S3087: begin
        IMAGE_addr <= 3071;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 732;
        test_state <= test_b1_S3088;
      end
      test_b1_S3088: begin
        IMAGE_addr <= 3072;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3089;
      end
      test_b1_S3089: begin
        IMAGE_addr <= 3073;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3090;
      end
      test_b1_S3090: begin
        IMAGE_addr <= 3074;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3047;
        test_state <= test_b1_S3091;
      end
      test_b1_S3091: begin
        IMAGE_addr <= 3075;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S3092;
      end
      test_b1_S3092: begin
        IMAGE_addr <= 3076;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3083;
        test_state <= test_b1_S3093;
      end
      test_b1_S3093: begin
        IMAGE_addr <= 3077;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 58;
        test_state <= test_b1_S3094;
      end
      test_b1_S3094: begin
        IMAGE_addr <= 3078;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 104;
        test_state <= test_b1_S3095;
      end
      test_b1_S3095: begin
        IMAGE_addr <= 3079;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S3096;
      end
      test_b1_S3096: begin
        IMAGE_addr <= 3080;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 100;
        test_state <= test_b1_S3097;
      end
      test_b1_S3097: begin
        IMAGE_addr <= 3081;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S3098;
      end
      test_b1_S3098: begin
        IMAGE_addr <= 3082;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3099;
      end
      test_b1_S3099: begin
        IMAGE_addr <= 3083;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3100;
      end
      test_b1_S3100: begin
        IMAGE_addr <= 3084;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3101;
      end
      test_b1_S3101: begin
        IMAGE_addr <= 3085;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S3102;
      end
      test_b1_S3102: begin
        IMAGE_addr <= 3086;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3056;
        test_state <= test_b1_S3103;
      end
      test_b1_S3103: begin
        IMAGE_addr <= 3087;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S3104;
      end
      test_b1_S3104: begin
        IMAGE_addr <= 3088;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S3105;
      end
      test_b1_S3105: begin
        IMAGE_addr <= 3089;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S3106;
      end
      test_b1_S3106: begin
        IMAGE_addr <= 3090;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 790;
        test_state <= test_b1_S3107;
      end
      test_b1_S3107: begin
        IMAGE_addr <= 3091;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S3108;
      end
      test_b1_S3108: begin
        IMAGE_addr <= 3092;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3102;
        test_state <= test_b1_S3109;
      end
      test_b1_S3109: begin
        IMAGE_addr <= 3093;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S3110;
      end
      test_b1_S3110: begin
        IMAGE_addr <= 3094;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S3111;
      end
      test_b1_S3111: begin
        IMAGE_addr <= 3095;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S3112;
      end
      test_b1_S3112: begin
        IMAGE_addr <= 3096;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S3113;
      end
      test_b1_S3113: begin
        IMAGE_addr <= 3097;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S3114;
      end
      test_b1_S3114: begin
        IMAGE_addr <= 3098;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S3115;
      end
      test_b1_S3115: begin
        IMAGE_addr <= 3099;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S3116;
      end
      test_b1_S3116: begin
        IMAGE_addr <= 3100;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S3117;
      end
      test_b1_S3117: begin
        IMAGE_addr <= 3101;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3118;
      end
      test_b1_S3118: begin
        IMAGE_addr <= 3102;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S3119;
      end
      test_b1_S3119: begin
        IMAGE_addr <= 3103;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3106;
        test_state <= test_b1_S3120;
      end
      test_b1_S3120: begin
        IMAGE_addr <= 3104;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3017;
        test_state <= test_b1_S3121;
      end
      test_b1_S3121: begin
        IMAGE_addr <= 3105;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3122;
      end
      test_b1_S3122: begin
        IMAGE_addr <= 3106;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 732;
        test_state <= test_b1_S3123;
      end
      test_b1_S3123: begin
        IMAGE_addr <= 3107;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3124;
      end
      test_b1_S3124: begin
        IMAGE_addr <= 3108;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3125;
      end
      test_b1_S3125: begin
        IMAGE_addr <= 3109;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3074;
        test_state <= test_b1_S3126;
      end
      test_b1_S3126: begin
        IMAGE_addr <= 3110;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S3127;
      end
      test_b1_S3127: begin
        IMAGE_addr <= 3111;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3117;
        test_state <= test_b1_S3128;
      end
      test_b1_S3128: begin
        IMAGE_addr <= 3112;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 104;
        test_state <= test_b1_S3129;
      end
      test_b1_S3129: begin
        IMAGE_addr <= 3113;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S3130;
      end
      test_b1_S3130: begin
        IMAGE_addr <= 3114;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 100;
        test_state <= test_b1_S3131;
      end
      test_b1_S3131: begin
        IMAGE_addr <= 3115;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S3132;
      end
      test_b1_S3132: begin
        IMAGE_addr <= 3116;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3133;
      end
      test_b1_S3133: begin
        IMAGE_addr <= 3117;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3134;
      end
      test_b1_S3134: begin
        IMAGE_addr <= 3118;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3135;
      end
      test_b1_S3135: begin
        IMAGE_addr <= 3119;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1239;
        test_state <= test_b1_S3136;
      end
      test_b1_S3136: begin
        IMAGE_addr <= 3120;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 25;
        test_state <= test_b1_S3137;
      end
      test_b1_S3137: begin
        IMAGE_addr <= 3121;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3083;
        test_state <= test_b1_S3138;
      end
      test_b1_S3138: begin
        IMAGE_addr <= 3122;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3139;
      end
      test_b1_S3139: begin
        IMAGE_addr <= 3123;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3140;
      end
      test_b1_S3140: begin
        IMAGE_addr <= 3124;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3109;
        test_state <= test_b1_S3141;
      end
      test_b1_S3141: begin
        IMAGE_addr <= 3125;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S3142;
      end
      test_b1_S3142: begin
        IMAGE_addr <= 3126;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3135;
        test_state <= test_b1_S3143;
      end
      test_b1_S3143: begin
        IMAGE_addr <= 3127;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S3144;
      end
      test_b1_S3144: begin
        IMAGE_addr <= 3128;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S3145;
      end
      test_b1_S3145: begin
        IMAGE_addr <= 3129;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 99;
        test_state <= test_b1_S3146;
      end
      test_b1_S3146: begin
        IMAGE_addr <= 3130;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 108;
        test_state <= test_b1_S3147;
      end
      test_b1_S3147: begin
        IMAGE_addr <= 3131;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S3148;
      end
      test_b1_S3148: begin
        IMAGE_addr <= 3132;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S3149;
      end
      test_b1_S3149: begin
        IMAGE_addr <= 3133;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S3150;
      end
      test_b1_S3150: begin
        IMAGE_addr <= 3134;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3151;
      end
      test_b1_S3151: begin
        IMAGE_addr <= 3135;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3152;
      end
      test_b1_S3152: begin
        IMAGE_addr <= 3136;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3153;
      end
      test_b1_S3153: begin
        IMAGE_addr <= 3137;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S3154;
      end
      test_b1_S3154: begin
        IMAGE_addr <= 3138;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S3155;
      end
      test_b1_S3155: begin
        IMAGE_addr <= 3139;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S3156;
      end
      test_b1_S3156: begin
        IMAGE_addr <= 3140;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 578;
        test_state <= test_b1_S3157;
      end
      test_b1_S3157: begin
        IMAGE_addr <= 3141;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S3158;
      end
      test_b1_S3158: begin
        IMAGE_addr <= 3142;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3159;
      end
      test_b1_S3159: begin
        IMAGE_addr <= 3143;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3160;
      end
      test_b1_S3160: begin
        IMAGE_addr <= 3144;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3124;
        test_state <= test_b1_S3161;
      end
      test_b1_S3161: begin
        IMAGE_addr <= 3145;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S3162;
      end
      test_b1_S3162: begin
        IMAGE_addr <= 3146;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3156;
        test_state <= test_b1_S3163;
      end
      test_b1_S3163: begin
        IMAGE_addr <= 3147;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S3164;
      end
      test_b1_S3164: begin
        IMAGE_addr <= 3148;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S3165;
      end
      test_b1_S3165: begin
        IMAGE_addr <= 3149;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 99;
        test_state <= test_b1_S3166;
      end
      test_b1_S3166: begin
        IMAGE_addr <= 3150;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 108;
        test_state <= test_b1_S3167;
      end
      test_b1_S3167: begin
        IMAGE_addr <= 3151;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S3168;
      end
      test_b1_S3168: begin
        IMAGE_addr <= 3152;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S3169;
      end
      test_b1_S3169: begin
        IMAGE_addr <= 3153;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S3170;
      end
      test_b1_S3170: begin
        IMAGE_addr <= 3154;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 58;
        test_state <= test_b1_S3171;
      end
      test_b1_S3171: begin
        IMAGE_addr <= 3155;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3172;
      end
      test_b1_S3172: begin
        IMAGE_addr <= 3156;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3173;
      end
      test_b1_S3173: begin
        IMAGE_addr <= 3157;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3174;
      end
      test_b1_S3174: begin
        IMAGE_addr <= 3158;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3038;
        test_state <= test_b1_S3175;
      end
      test_b1_S3175: begin
        IMAGE_addr <= 3159;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 578;
        test_state <= test_b1_S3176;
      end
      test_b1_S3176: begin
        IMAGE_addr <= 3160;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S3177;
      end
      test_b1_S3177: begin
        IMAGE_addr <= 3161;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3178;
      end
      test_b1_S3178: begin
        IMAGE_addr <= 3162;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3179;
      end
      test_b1_S3179: begin
        IMAGE_addr <= 3163;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3144;
        test_state <= test_b1_S3180;
      end
      test_b1_S3180: begin
        IMAGE_addr <= 3164;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S3181;
      end
      test_b1_S3181: begin
        IMAGE_addr <= 3165;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3175;
        test_state <= test_b1_S3182;
      end
      test_b1_S3182: begin
        IMAGE_addr <= 3166;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 120;
        test_state <= test_b1_S3183;
      end
      test_b1_S3183: begin
        IMAGE_addr <= 3167;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S3184;
      end
      test_b1_S3184: begin
        IMAGE_addr <= 3168;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 58;
        test_state <= test_b1_S3185;
      end
      test_b1_S3185: begin
        IMAGE_addr <= 3169;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 99;
        test_state <= test_b1_S3186;
      end
      test_b1_S3186: begin
        IMAGE_addr <= 3170;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 108;
        test_state <= test_b1_S3187;
      end
      test_b1_S3187: begin
        IMAGE_addr <= 3171;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S3188;
      end
      test_b1_S3188: begin
        IMAGE_addr <= 3172;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S3189;
      end
      test_b1_S3189: begin
        IMAGE_addr <= 3173;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S3190;
      end
      test_b1_S3190: begin
        IMAGE_addr <= 3174;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3191;
      end
      test_b1_S3191: begin
        IMAGE_addr <= 3175;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S3192;
      end
      test_b1_S3192: begin
        IMAGE_addr <= 3176;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3056;
        test_state <= test_b1_S3193;
      end
      test_b1_S3193: begin
        IMAGE_addr <= 3177;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 25;
        test_state <= test_b1_S3194;
      end
      test_b1_S3194: begin
        IMAGE_addr <= 3178;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 578;
        test_state <= test_b1_S3195;
      end
      test_b1_S3195: begin
        IMAGE_addr <= 3179;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S3196;
      end
      test_b1_S3196: begin
        IMAGE_addr <= 3180;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 286;
        test_state <= test_b1_S3197;
      end
      test_b1_S3197: begin
        IMAGE_addr <= 3181;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3198;
      end
      test_b1_S3198: begin
        IMAGE_addr <= 3182;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3199;
      end
      test_b1_S3199: begin
        IMAGE_addr <= 3183;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3144;
        test_state <= test_b1_S3200;
      end
      test_b1_S3200: begin
        IMAGE_addr <= 3184;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 306;
        test_state <= test_b1_S3201;
      end
      test_b1_S3201: begin
        IMAGE_addr <= 3185;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3190;
        test_state <= test_b1_S3202;
      end
      test_b1_S3202: begin
        IMAGE_addr <= 3186;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 95;
        test_state <= test_b1_S3203;
      end
      test_b1_S3203: begin
        IMAGE_addr <= 3187;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 95;
        test_state <= test_b1_S3204;
      end
      test_b1_S3204: begin
        IMAGE_addr <= 3188;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 38;
        test_state <= test_b1_S3205;
      end
      test_b1_S3205: begin
        IMAGE_addr <= 3189;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3206;
      end
      test_b1_S3206: begin
        IMAGE_addr <= 3190;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3207;
      end
      test_b1_S3207: begin
        IMAGE_addr <= 3191;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3208;
      end
      test_b1_S3208: begin
        IMAGE_addr <= 3192;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 310;
        test_state <= test_b1_S3209;
      end
      test_b1_S3209: begin
        IMAGE_addr <= 3193;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3210;
      end
      test_b1_S3210: begin
        IMAGE_addr <= 3194;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3211;
      end
      test_b1_S3211: begin
        IMAGE_addr <= 3195;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3183;
        test_state <= test_b1_S3212;
      end
      test_b1_S3212: begin
        IMAGE_addr <= 3196;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 306;
        test_state <= test_b1_S3213;
      end
      test_b1_S3213: begin
        IMAGE_addr <= 3197;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3202;
        test_state <= test_b1_S3214;
      end
      test_b1_S3214: begin
        IMAGE_addr <= 3198;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 95;
        test_state <= test_b1_S3215;
      end
      test_b1_S3215: begin
        IMAGE_addr <= 3199;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 95;
        test_state <= test_b1_S3216;
      end
      test_b1_S3216: begin
        IMAGE_addr <= 3200;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 64;
        test_state <= test_b1_S3217;
      end
      test_b1_S3217: begin
        IMAGE_addr <= 3201;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3218;
      end
      test_b1_S3218: begin
        IMAGE_addr <= 3202;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3219;
      end
      test_b1_S3219: begin
        IMAGE_addr <= 3203;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3220;
      end
      test_b1_S3220: begin
        IMAGE_addr <= 3204;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3175;
        test_state <= test_b1_S3221;
      end
      test_b1_S3221: begin
        IMAGE_addr <= 3205;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S3222;
      end
      test_b1_S3222: begin
        IMAGE_addr <= 3206;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 72;
        test_state <= test_b1_S3223;
      end
      test_b1_S3223: begin
        IMAGE_addr <= 3207;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3175;
        test_state <= test_b1_S3224;
      end
      test_b1_S3224: begin
        IMAGE_addr <= 3208;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3225;
      end
      test_b1_S3225: begin
        IMAGE_addr <= 3209;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3226;
      end
      test_b1_S3226: begin
        IMAGE_addr <= 3210;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3195;
        test_state <= test_b1_S3227;
      end
      test_b1_S3227: begin
        IMAGE_addr <= 3211;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 306;
        test_state <= test_b1_S3228;
      end
      test_b1_S3228: begin
        IMAGE_addr <= 3212;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3217;
        test_state <= test_b1_S3229;
      end
      test_b1_S3229: begin
        IMAGE_addr <= 3213;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 95;
        test_state <= test_b1_S3230;
      end
      test_b1_S3230: begin
        IMAGE_addr <= 3214;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 95;
        test_state <= test_b1_S3231;
      end
      test_b1_S3231: begin
        IMAGE_addr <= 3215;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 33;
        test_state <= test_b1_S3232;
      end
      test_b1_S3232: begin
        IMAGE_addr <= 3216;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3233;
      end
      test_b1_S3233: begin
        IMAGE_addr <= 3217;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3234;
      end
      test_b1_S3234: begin
        IMAGE_addr <= 3218;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3235;
      end
      test_b1_S3235: begin
        IMAGE_addr <= 3219;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3175;
        test_state <= test_b1_S3236;
      end
      test_b1_S3236: begin
        IMAGE_addr <= 3220;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S3237;
      end
      test_b1_S3237: begin
        IMAGE_addr <= 3221;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 77;
        test_state <= test_b1_S3238;
      end
      test_b1_S3238: begin
        IMAGE_addr <= 3222;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3175;
        test_state <= test_b1_S3239;
      end
      test_b1_S3239: begin
        IMAGE_addr <= 3223;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3240;
      end
      test_b1_S3240: begin
        IMAGE_addr <= 3224;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3241;
      end
      test_b1_S3241: begin
        IMAGE_addr <= 3225;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3210;
        test_state <= test_b1_S3242;
      end
      test_b1_S3242: begin
        IMAGE_addr <= 3226;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 306;
        test_state <= test_b1_S3243;
      end
      test_b1_S3243: begin
        IMAGE_addr <= 3227;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3232;
        test_state <= test_b1_S3244;
      end
      test_b1_S3244: begin
        IMAGE_addr <= 3228;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 95;
        test_state <= test_b1_S3245;
      end
      test_b1_S3245: begin
        IMAGE_addr <= 3229;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 95;
        test_state <= test_b1_S3246;
      end
      test_b1_S3246: begin
        IMAGE_addr <= 3230;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 43;
        test_state <= test_b1_S3247;
      end
      test_b1_S3247: begin
        IMAGE_addr <= 3231;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3248;
      end
      test_b1_S3248: begin
        IMAGE_addr <= 3232;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3249;
      end
      test_b1_S3249: begin
        IMAGE_addr <= 3233;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3250;
      end
      test_b1_S3250: begin
        IMAGE_addr <= 3234;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3175;
        test_state <= test_b1_S3251;
      end
      test_b1_S3251: begin
        IMAGE_addr <= 3235;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S3252;
      end
      test_b1_S3252: begin
        IMAGE_addr <= 3236;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2618;
        test_state <= test_b1_S3253;
      end
      test_b1_S3253: begin
        IMAGE_addr <= 3237;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S3254;
      end
      test_b1_S3254: begin
        IMAGE_addr <= 3238;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3255;
      end
      test_b1_S3255: begin
        IMAGE_addr <= 3239;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3256;
      end
      test_b1_S3256: begin
        IMAGE_addr <= 3240;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3225;
        test_state <= test_b1_S3257;
      end
      test_b1_S3257: begin
        IMAGE_addr <= 3241;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 306;
        test_state <= test_b1_S3258;
      end
      test_b1_S3258: begin
        IMAGE_addr <= 3242;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3247;
        test_state <= test_b1_S3259;
      end
      test_b1_S3259: begin
        IMAGE_addr <= 3243;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 95;
        test_state <= test_b1_S3260;
      end
      test_b1_S3260: begin
        IMAGE_addr <= 3244;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 95;
        test_state <= test_b1_S3261;
      end
      test_b1_S3261: begin
        IMAGE_addr <= 3245;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 45;
        test_state <= test_b1_S3262;
      end
      test_b1_S3262: begin
        IMAGE_addr <= 3246;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3263;
      end
      test_b1_S3263: begin
        IMAGE_addr <= 3247;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3264;
      end
      test_b1_S3264: begin
        IMAGE_addr <= 3248;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3265;
      end
      test_b1_S3265: begin
        IMAGE_addr <= 3249;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3175;
        test_state <= test_b1_S3266;
      end
      test_b1_S3266: begin
        IMAGE_addr <= 3250;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S3267;
      end
      test_b1_S3267: begin
        IMAGE_addr <= 3251;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2634;
        test_state <= test_b1_S3268;
      end
      test_b1_S3268: begin
        IMAGE_addr <= 3252;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S3269;
      end
      test_b1_S3269: begin
        IMAGE_addr <= 3253;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3270;
      end
      test_b1_S3270: begin
        IMAGE_addr <= 3254;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3271;
      end
      test_b1_S3271: begin
        IMAGE_addr <= 3255;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3240;
        test_state <= test_b1_S3272;
      end
      test_b1_S3272: begin
        IMAGE_addr <= 3256;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 306;
        test_state <= test_b1_S3273;
      end
      test_b1_S3273: begin
        IMAGE_addr <= 3257;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3262;
        test_state <= test_b1_S3274;
      end
      test_b1_S3274: begin
        IMAGE_addr <= 3258;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 95;
        test_state <= test_b1_S3275;
      end
      test_b1_S3275: begin
        IMAGE_addr <= 3259;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 95;
        test_state <= test_b1_S3276;
      end
      test_b1_S3276: begin
        IMAGE_addr <= 3260;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 50;
        test_state <= test_b1_S3277;
      end
      test_b1_S3277: begin
        IMAGE_addr <= 3261;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3278;
      end
      test_b1_S3278: begin
        IMAGE_addr <= 3262;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3279;
      end
      test_b1_S3279: begin
        IMAGE_addr <= 3263;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3280;
      end
      test_b1_S3280: begin
        IMAGE_addr <= 3264;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S3281;
      end
      test_b1_S3281: begin
        IMAGE_addr <= 3265;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3175;
        test_state <= test_b1_S3282;
      end
      test_b1_S3282: begin
        IMAGE_addr <= 3266;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 774;
        test_state <= test_b1_S3283;
      end
      test_b1_S3283: begin
        IMAGE_addr <= 3267;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3175;
        test_state <= test_b1_S3284;
      end
      test_b1_S3284: begin
        IMAGE_addr <= 3268;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3285;
      end
      test_b1_S3285: begin
        IMAGE_addr <= 3269;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3286;
      end
      test_b1_S3286: begin
        IMAGE_addr <= 3270;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3255;
        test_state <= test_b1_S3287;
      end
      test_b1_S3287: begin
        IMAGE_addr <= 3271;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S3288;
      end
      test_b1_S3288: begin
        IMAGE_addr <= 3272;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3283;
        test_state <= test_b1_S3289;
      end
      test_b1_S3289: begin
        IMAGE_addr <= 3273;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 46;
        test_state <= test_b1_S3290;
      end
      test_b1_S3290: begin
        IMAGE_addr <= 3274;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 99;
        test_state <= test_b1_S3291;
      end
      test_b1_S3291: begin
        IMAGE_addr <= 3275;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 111;
        test_state <= test_b1_S3292;
      end
      test_b1_S3292: begin
        IMAGE_addr <= 3276;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 109;
        test_state <= test_b1_S3293;
      end
      test_b1_S3293: begin
        IMAGE_addr <= 3277;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 112;
        test_state <= test_b1_S3294;
      end
      test_b1_S3294: begin
        IMAGE_addr <= 3278;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S3295;
      end
      test_b1_S3295: begin
        IMAGE_addr <= 3279;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 108;
        test_state <= test_b1_S3296;
      end
      test_b1_S3296: begin
        IMAGE_addr <= 3280;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S3297;
      end
      test_b1_S3297: begin
        IMAGE_addr <= 3281;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S3298;
      end
      test_b1_S3298: begin
        IMAGE_addr <= 3282;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3299;
      end
      test_b1_S3299: begin
        IMAGE_addr <= 3283;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3300;
      end
      test_b1_S3300: begin
        IMAGE_addr <= 3284;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3301;
      end
      test_b1_S3301: begin
        IMAGE_addr <= 3285;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S3302;
      end
      test_b1_S3302: begin
        IMAGE_addr <= 3286;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S3303;
      end
      test_b1_S3303: begin
        IMAGE_addr <= 3287;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S3304;
      end
      test_b1_S3304: begin
        IMAGE_addr <= 3288;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S3305;
      end
      test_b1_S3305: begin
        IMAGE_addr <= 3289;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 183;
        test_state <= test_b1_S3306;
      end
      test_b1_S3306: begin
        IMAGE_addr <= 3290;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S3307;
      end
      test_b1_S3307: begin
        IMAGE_addr <= 3291;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 52;
        test_state <= test_b1_S3308;
      end
      test_b1_S3308: begin
        IMAGE_addr <= 3292;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 732;
        test_state <= test_b1_S3309;
      end
      test_b1_S3309: begin
        IMAGE_addr <= 3293;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3310;
      end
      test_b1_S3310: begin
        IMAGE_addr <= 3294;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3311;
      end
      test_b1_S3311: begin
        IMAGE_addr <= 3295;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3270;
        test_state <= test_b1_S3312;
      end
      test_b1_S3312: begin
        IMAGE_addr <= 3296;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S3313;
      end
      test_b1_S3313: begin
        IMAGE_addr <= 3297;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3308;
        test_state <= test_b1_S3314;
      end
      test_b1_S3314: begin
        IMAGE_addr <= 3298;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S3315;
      end
      test_b1_S3315: begin
        IMAGE_addr <= 3299;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 109;
        test_state <= test_b1_S3316;
      end
      test_b1_S3316: begin
        IMAGE_addr <= 3300;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 109;
        test_state <= test_b1_S3317;
      end
      test_b1_S3317: begin
        IMAGE_addr <= 3301;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S3318;
      end
      test_b1_S3318: begin
        IMAGE_addr <= 3302;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 100;
        test_state <= test_b1_S3319;
      end
      test_b1_S3319: begin
        IMAGE_addr <= 3303;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S3320;
      end
      test_b1_S3320: begin
        IMAGE_addr <= 3304;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S3321;
      end
      test_b1_S3321: begin
        IMAGE_addr <= 3305;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S3322;
      end
      test_b1_S3322: begin
        IMAGE_addr <= 3306;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S3323;
      end
      test_b1_S3323: begin
        IMAGE_addr <= 3307;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3324;
      end
      test_b1_S3324: begin
        IMAGE_addr <= 3308;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3325;
      end
      test_b1_S3325: begin
        IMAGE_addr <= 3309;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3326;
      end
      test_b1_S3326: begin
        IMAGE_addr <= 3310;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S3327;
      end
      test_b1_S3327: begin
        IMAGE_addr <= 3311;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 306;
        test_state <= test_b1_S3328;
      end
      test_b1_S3328: begin
        IMAGE_addr <= 3312;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3135;
        test_state <= test_b1_S3329;
      end
      test_b1_S3329: begin
        IMAGE_addr <= 3313;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3330;
      end
      test_b1_S3330: begin
        IMAGE_addr <= 3314;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3331;
      end
      test_b1_S3331: begin
        IMAGE_addr <= 3315;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3295;
        test_state <= test_b1_S3332;
      end
      test_b1_S3332: begin
        IMAGE_addr <= 3316;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S3333;
      end
      test_b1_S3333: begin
        IMAGE_addr <= 3317;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3331;
        test_state <= test_b1_S3334;
      end
      test_b1_S3334: begin
        IMAGE_addr <= 3318;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 99;
        test_state <= test_b1_S3335;
      end
      test_b1_S3335: begin
        IMAGE_addr <= 3319;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 111;
        test_state <= test_b1_S3336;
      end
      test_b1_S3336: begin
        IMAGE_addr <= 3320;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 109;
        test_state <= test_b1_S3337;
      end
      test_b1_S3337: begin
        IMAGE_addr <= 3321;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 112;
        test_state <= test_b1_S3338;
      end
      test_b1_S3338: begin
        IMAGE_addr <= 3322;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S3339;
      end
      test_b1_S3339: begin
        IMAGE_addr <= 3323;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 108;
        test_state <= test_b1_S3340;
      end
      test_b1_S3340: begin
        IMAGE_addr <= 3324;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S3341;
      end
      test_b1_S3341: begin
        IMAGE_addr <= 3325;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 45;
        test_state <= test_b1_S3342;
      end
      test_b1_S3342: begin
        IMAGE_addr <= 3326;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 111;
        test_state <= test_b1_S3343;
      end
      test_b1_S3343: begin
        IMAGE_addr <= 3327;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 110;
        test_state <= test_b1_S3344;
      end
      test_b1_S3344: begin
        IMAGE_addr <= 3328;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 108;
        test_state <= test_b1_S3345;
      end
      test_b1_S3345: begin
        IMAGE_addr <= 3329;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 121;
        test_state <= test_b1_S3346;
      end
      test_b1_S3346: begin
        IMAGE_addr <= 3330;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3347;
      end
      test_b1_S3347: begin
        IMAGE_addr <= 3331;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3348;
      end
      test_b1_S3348: begin
        IMAGE_addr <= 3332;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3349;
      end
      test_b1_S3349: begin
        IMAGE_addr <= 3333;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S3350;
      end
      test_b1_S3350: begin
        IMAGE_addr <= 3334;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3283;
        test_state <= test_b1_S3351;
      end
      test_b1_S3351: begin
        IMAGE_addr <= 3335;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3135;
        test_state <= test_b1_S3352;
      end
      test_b1_S3352: begin
        IMAGE_addr <= 3336;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3353;
      end
      test_b1_S3353: begin
        IMAGE_addr <= 3337;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3354;
      end
      test_b1_S3354: begin
        IMAGE_addr <= 3338;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3315;
        test_state <= test_b1_S3355;
      end
      test_b1_S3355: begin
        IMAGE_addr <= 3339;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3283;
        test_state <= test_b1_S3356;
      end
      test_b1_S3356: begin
        IMAGE_addr <= 3340;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3343;
        test_state <= test_b1_S3357;
      end
      test_b1_S3357: begin
        IMAGE_addr <= 3341;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 96;
        test_state <= test_b1_S3358;
      end
      test_b1_S3358: begin
        IMAGE_addr <= 3342;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3359;
      end
      test_b1_S3359: begin
        IMAGE_addr <= 3343;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3360;
      end
      test_b1_S3360: begin
        IMAGE_addr <= 3344;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3361;
      end
      test_b1_S3361: begin
        IMAGE_addr <= 3345;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1239;
        test_state <= test_b1_S3362;
      end
      test_b1_S3362: begin
        IMAGE_addr <= 3346;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S3363;
      end
      test_b1_S3363: begin
        IMAGE_addr <= 3347;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S3364;
      end
      test_b1_S3364: begin
        IMAGE_addr <= 3348;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3365;
      end
      test_b1_S3365: begin
        IMAGE_addr <= 3349;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 798;
        test_state <= test_b1_S3366;
      end
      test_b1_S3366: begin
        IMAGE_addr <= 3350;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S3367;
      end
      test_b1_S3367: begin
        IMAGE_addr <= 3351;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4294967295;
        test_state <= test_b1_S3368;
      end
      test_b1_S3368: begin
        IMAGE_addr <= 3352;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 790;
        test_state <= test_b1_S3369;
      end
      test_b1_S3369: begin
        IMAGE_addr <= 3353;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S3370;
      end
      test_b1_S3370: begin
        IMAGE_addr <= 3354;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3363;
        test_state <= test_b1_S3371;
      end
      test_b1_S3371: begin
        IMAGE_addr <= 3355;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 310;
        test_state <= test_b1_S3372;
      end
      test_b1_S3372: begin
        IMAGE_addr <= 3356;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S3373;
      end
      test_b1_S3373: begin
        IMAGE_addr <= 3357;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5;
        test_state <= test_b1_S3374;
      end
      test_b1_S3374: begin
        IMAGE_addr <= 3358;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S3375;
      end
      test_b1_S3375: begin
        IMAGE_addr <= 3359;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 578;
        test_state <= test_b1_S3376;
      end
      test_b1_S3376: begin
        IMAGE_addr <= 3360;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S3377;
      end
      test_b1_S3377: begin
        IMAGE_addr <= 3361;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 213;
        test_state <= test_b1_S3378;
      end
      test_b1_S3378: begin
        IMAGE_addr <= 3362;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3379;
      end
      test_b1_S3379: begin
        IMAGE_addr <= 3363;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S3380;
      end
      test_b1_S3380: begin
        IMAGE_addr <= 3364;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3386;
        test_state <= test_b1_S3381;
      end
      test_b1_S3381: begin
        IMAGE_addr <= 3365;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S3382;
      end
      test_b1_S3382: begin
        IMAGE_addr <= 3366;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 400;
        test_state <= test_b1_S3383;
      end
      test_b1_S3383: begin
        IMAGE_addr <= 3367;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1091;
        test_state <= test_b1_S3384;
      end
      test_b1_S3384: begin
        IMAGE_addr <= 3368;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S3385;
      end
      test_b1_S3385: begin
        IMAGE_addr <= 3369;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4294967295;
        test_state <= test_b1_S3386;
      end
      test_b1_S3386: begin
        IMAGE_addr <= 3370;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 790;
        test_state <= test_b1_S3387;
      end
      test_b1_S3387: begin
        IMAGE_addr <= 3371;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S3388;
      end
      test_b1_S3388: begin
        IMAGE_addr <= 3372;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3380;
        test_state <= test_b1_S3389;
      end
      test_b1_S3389: begin
        IMAGE_addr <= 3373;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 400;
        test_state <= test_b1_S3390;
      end
      test_b1_S3390: begin
        IMAGE_addr <= 3374;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1056;
        test_state <= test_b1_S3391;
      end
      test_b1_S3391: begin
        IMAGE_addr <= 3375;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 310;
        test_state <= test_b1_S3392;
      end
      test_b1_S3392: begin
        IMAGE_addr <= 3376;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S3393;
      end
      test_b1_S3393: begin
        IMAGE_addr <= 3377;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 310;
        test_state <= test_b1_S3394;
      end
      test_b1_S3394: begin
        IMAGE_addr <= 3378;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 213;
        test_state <= test_b1_S3395;
      end
      test_b1_S3395: begin
        IMAGE_addr <= 3379;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3396;
      end
      test_b1_S3396: begin
        IMAGE_addr <= 3380;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S3397;
      end
      test_b1_S3397: begin
        IMAGE_addr <= 3381;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3384;
        test_state <= test_b1_S3398;
      end
      test_b1_S3398: begin
        IMAGE_addr <= 3382;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1321;
        test_state <= test_b1_S3399;
      end
      test_b1_S3399: begin
        IMAGE_addr <= 3383;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3400;
      end
      test_b1_S3400: begin
        IMAGE_addr <= 3384;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 732;
        test_state <= test_b1_S3401;
      end
      test_b1_S3401: begin
        IMAGE_addr <= 3385;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3402;
      end
      test_b1_S3402: begin
        IMAGE_addr <= 3386;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 732;
        test_state <= test_b1_S3403;
      end
      test_b1_S3403: begin
        IMAGE_addr <= 3387;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3404;
      end
      test_b1_S3404: begin
        IMAGE_addr <= 3388;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3405;
      end
      test_b1_S3405: begin
        IMAGE_addr <= 3389;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3338;
        test_state <= test_b1_S3406;
      end
      test_b1_S3406: begin
        IMAGE_addr <= 3390;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3283;
        test_state <= test_b1_S3407;
      end
      test_b1_S3407: begin
        IMAGE_addr <= 3391;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3398;
        test_state <= test_b1_S3408;
      end
      test_b1_S3408: begin
        IMAGE_addr <= 3392;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 106;
        test_state <= test_b1_S3409;
      end
      test_b1_S3409: begin
        IMAGE_addr <= 3393;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 117;
        test_state <= test_b1_S3410;
      end
      test_b1_S3410: begin
        IMAGE_addr <= 3394;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 109;
        test_state <= test_b1_S3411;
      end
      test_b1_S3411: begin
        IMAGE_addr <= 3395;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 112;
        test_state <= test_b1_S3412;
      end
      test_b1_S3412: begin
        IMAGE_addr <= 3396;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 58;
        test_state <= test_b1_S3413;
      end
      test_b1_S3413: begin
        IMAGE_addr <= 3397;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3414;
      end
      test_b1_S3414: begin
        IMAGE_addr <= 3398;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3415;
      end
      test_b1_S3415: begin
        IMAGE_addr <= 3399;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3416;
      end
      test_b1_S3416: begin
        IMAGE_addr <= 3400;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1239;
        test_state <= test_b1_S3417;
      end
      test_b1_S3417: begin
        IMAGE_addr <= 3401;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 25;
        test_state <= test_b1_S3418;
      end
      test_b1_S3418: begin
        IMAGE_addr <= 3402;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S3419;
      end
      test_b1_S3419: begin
        IMAGE_addr <= 3403;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8;
        test_state <= test_b1_S3420;
      end
      test_b1_S3420: begin
        IMAGE_addr <= 3404;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 213;
        test_state <= test_b1_S3421;
      end
      test_b1_S3421: begin
        IMAGE_addr <= 3405;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 213;
        test_state <= test_b1_S3422;
      end
      test_b1_S3422: begin
        IMAGE_addr <= 3406;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3423;
      end
      test_b1_S3423: begin
        IMAGE_addr <= 3407;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3424;
      end
      test_b1_S3424: begin
        IMAGE_addr <= 3408;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3389;
        test_state <= test_b1_S3425;
      end
      test_b1_S3425: begin
        IMAGE_addr <= 3409;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 306;
        test_state <= test_b1_S3426;
      end
      test_b1_S3426: begin
        IMAGE_addr <= 3410;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3414;
        test_state <= test_b1_S3427;
      end
      test_b1_S3427: begin
        IMAGE_addr <= 3411;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 91;
        test_state <= test_b1_S3428;
      end
      test_b1_S3428: begin
        IMAGE_addr <= 3412;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 93;
        test_state <= test_b1_S3429;
      end
      test_b1_S3429: begin
        IMAGE_addr <= 3413;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3430;
      end
      test_b1_S3430: begin
        IMAGE_addr <= 3414;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3431;
      end
      test_b1_S3431: begin
        IMAGE_addr <= 3415;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3432;
      end
      test_b1_S3432: begin
        IMAGE_addr <= 3416;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S3433;
      end
      test_b1_S3433: begin
        IMAGE_addr <= 3417;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 691;
        test_state <= test_b1_S3434;
      end
      test_b1_S3434: begin
        IMAGE_addr <= 3418;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 306;
        test_state <= test_b1_S3435;
      end
      test_b1_S3435: begin
        IMAGE_addr <= 3419;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S3436;
      end
      test_b1_S3436: begin
        IMAGE_addr <= 3420;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 708;
        test_state <= test_b1_S3437;
      end
      test_b1_S3437: begin
        IMAGE_addr <= 3421;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 306;
        test_state <= test_b1_S3438;
      end
      test_b1_S3438: begin
        IMAGE_addr <= 3422;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3439;
      end
      test_b1_S3439: begin
        IMAGE_addr <= 3423;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3440;
      end
      test_b1_S3440: begin
        IMAGE_addr <= 3424;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3408;
        test_state <= test_b1_S3441;
      end
      test_b1_S3441: begin
        IMAGE_addr <= 3425;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S3442;
      end
      test_b1_S3442: begin
        IMAGE_addr <= 3426;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3433;
        test_state <= test_b1_S3443;
      end
      test_b1_S3443: begin
        IMAGE_addr <= 3427;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 119;
        test_state <= test_b1_S3444;
      end
      test_b1_S3444: begin
        IMAGE_addr <= 3428;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 104;
        test_state <= test_b1_S3445;
      end
      test_b1_S3445: begin
        IMAGE_addr <= 3429;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S3446;
      end
      test_b1_S3446: begin
        IMAGE_addr <= 3430;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 108;
        test_state <= test_b1_S3447;
      end
      test_b1_S3447: begin
        IMAGE_addr <= 3431;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S3448;
      end
      test_b1_S3448: begin
        IMAGE_addr <= 3432;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3449;
      end
      test_b1_S3449: begin
        IMAGE_addr <= 3433;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3450;
      end
      test_b1_S3450: begin
        IMAGE_addr <= 3434;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3451;
      end
      test_b1_S3451: begin
        IMAGE_addr <= 3435;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S3452;
      end
      test_b1_S3452: begin
        IMAGE_addr <= 3436;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3445;
        test_state <= test_b1_S3453;
      end
      test_b1_S3453: begin
        IMAGE_addr <= 3437;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S3454;
      end
      test_b1_S3454: begin
        IMAGE_addr <= 3438;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 766;
        test_state <= test_b1_S3455;
      end
      test_b1_S3455: begin
        IMAGE_addr <= 3439;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S3456;
      end
      test_b1_S3456: begin
        IMAGE_addr <= 3440;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 25;
        test_state <= test_b1_S3457;
      end
      test_b1_S3457: begin
        IMAGE_addr <= 3441;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S3458;
      end
      test_b1_S3458: begin
        IMAGE_addr <= 3442;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8;
        test_state <= test_b1_S3459;
      end
      test_b1_S3459: begin
        IMAGE_addr <= 3443;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3437;
        test_state <= test_b1_S3460;
      end
      test_b1_S3460: begin
        IMAGE_addr <= 3444;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3461;
      end
      test_b1_S3461: begin
        IMAGE_addr <= 3445;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 183;
        test_state <= test_b1_S3462;
      end
      test_b1_S3462: begin
        IMAGE_addr <= 3446;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S3463;
      end
      test_b1_S3463: begin
        IMAGE_addr <= 3447;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3464;
      end
      test_b1_S3464: begin
        IMAGE_addr <= 3448;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3465;
      end
      test_b1_S3465: begin
        IMAGE_addr <= 3449;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3424;
        test_state <= test_b1_S3466;
      end
      test_b1_S3466: begin
        IMAGE_addr <= 3450;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S3467;
      end
      test_b1_S3467: begin
        IMAGE_addr <= 3451;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3458;
        test_state <= test_b1_S3468;
      end
      test_b1_S3468: begin
        IMAGE_addr <= 3452;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 117;
        test_state <= test_b1_S3469;
      end
      test_b1_S3469: begin
        IMAGE_addr <= 3453;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 110;
        test_state <= test_b1_S3470;
      end
      test_b1_S3470: begin
        IMAGE_addr <= 3454;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S3471;
      end
      test_b1_S3471: begin
        IMAGE_addr <= 3455;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S3472;
      end
      test_b1_S3472: begin
        IMAGE_addr <= 3456;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 108;
        test_state <= test_b1_S3473;
      end
      test_b1_S3473: begin
        IMAGE_addr <= 3457;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3474;
      end
      test_b1_S3474: begin
        IMAGE_addr <= 3458;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3475;
      end
      test_b1_S3475: begin
        IMAGE_addr <= 3459;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3476;
      end
      test_b1_S3476: begin
        IMAGE_addr <= 3460;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S3477;
      end
      test_b1_S3477: begin
        IMAGE_addr <= 3461;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3471;
        test_state <= test_b1_S3478;
      end
      test_b1_S3478: begin
        IMAGE_addr <= 3462;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S3479;
      end
      test_b1_S3479: begin
        IMAGE_addr <= 3463;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 766;
        test_state <= test_b1_S3480;
      end
      test_b1_S3480: begin
        IMAGE_addr <= 3464;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S3481;
      end
      test_b1_S3481: begin
        IMAGE_addr <= 3465;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 140;
        test_state <= test_b1_S3482;
      end
      test_b1_S3482: begin
        IMAGE_addr <= 3466;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 25;
        test_state <= test_b1_S3483;
      end
      test_b1_S3483: begin
        IMAGE_addr <= 3467;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S3484;
      end
      test_b1_S3484: begin
        IMAGE_addr <= 3468;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8;
        test_state <= test_b1_S3485;
      end
      test_b1_S3485: begin
        IMAGE_addr <= 3469;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3462;
        test_state <= test_b1_S3486;
      end
      test_b1_S3486: begin
        IMAGE_addr <= 3470;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3487;
      end
      test_b1_S3487: begin
        IMAGE_addr <= 3471;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 183;
        test_state <= test_b1_S3488;
      end
      test_b1_S3488: begin
        IMAGE_addr <= 3472;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S3489;
      end
      test_b1_S3489: begin
        IMAGE_addr <= 3473;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3490;
      end
      test_b1_S3490: begin
        IMAGE_addr <= 3474;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3491;
      end
      test_b1_S3491: begin
        IMAGE_addr <= 3475;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3449;
        test_state <= test_b1_S3492;
      end
      test_b1_S3492: begin
        IMAGE_addr <= 3476;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S3493;
      end
      test_b1_S3493: begin
        IMAGE_addr <= 3477;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3484;
        test_state <= test_b1_S3494;
      end
      test_b1_S3494: begin
        IMAGE_addr <= 3478;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 99;
        test_state <= test_b1_S3495;
      end
      test_b1_S3495: begin
        IMAGE_addr <= 3479;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 117;
        test_state <= test_b1_S3496;
      end
      test_b1_S3496: begin
        IMAGE_addr <= 3480;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S3497;
      end
      test_b1_S3497: begin
        IMAGE_addr <= 3481;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S3498;
      end
      test_b1_S3498: begin
        IMAGE_addr <= 3482;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 121;
        test_state <= test_b1_S3499;
      end
      test_b1_S3499: begin
        IMAGE_addr <= 3483;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3500;
      end
      test_b1_S3500: begin
        IMAGE_addr <= 3484;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3501;
      end
      test_b1_S3501: begin
        IMAGE_addr <= 3485;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3502;
      end
      test_b1_S3502: begin
        IMAGE_addr <= 3486;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S3503;
      end
      test_b1_S3503: begin
        IMAGE_addr <= 3487;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3497;
        test_state <= test_b1_S3504;
      end
      test_b1_S3504: begin
        IMAGE_addr <= 3488;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S3505;
      end
      test_b1_S3505: begin
        IMAGE_addr <= 3489;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3494;
        test_state <= test_b1_S3506;
      end
      test_b1_S3506: begin
        IMAGE_addr <= 3490;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S3507;
      end
      test_b1_S3507: begin
        IMAGE_addr <= 3491;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 691;
        test_state <= test_b1_S3508;
      end
      test_b1_S3508: begin
        IMAGE_addr <= 3492;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 306;
        test_state <= test_b1_S3509;
      end
      test_b1_S3509: begin
        IMAGE_addr <= 3493;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3510;
      end
      test_b1_S3510: begin
        IMAGE_addr <= 3494;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 766;
        test_state <= test_b1_S3511;
      end
      test_b1_S3511: begin
        IMAGE_addr <= 3495;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 310;
        test_state <= test_b1_S3512;
      end
      test_b1_S3512: begin
        IMAGE_addr <= 3496;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3513;
      end
      test_b1_S3513: begin
        IMAGE_addr <= 3497;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 766;
        test_state <= test_b1_S3514;
      end
      test_b1_S3514: begin
        IMAGE_addr <= 3498;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 213;
        test_state <= test_b1_S3515;
      end
      test_b1_S3515: begin
        IMAGE_addr <= 3499;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S3516;
      end
      test_b1_S3516: begin
        IMAGE_addr <= 3500;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 708;
        test_state <= test_b1_S3517;
      end
      test_b1_S3517: begin
        IMAGE_addr <= 3501;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 306;
        test_state <= test_b1_S3518;
      end
      test_b1_S3518: begin
        IMAGE_addr <= 3502;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3519;
      end
      test_b1_S3519: begin
        IMAGE_addr <= 3503;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3520;
      end
      test_b1_S3520: begin
        IMAGE_addr <= 3504;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3475;
        test_state <= test_b1_S3521;
      end
      test_b1_S3521: begin
        IMAGE_addr <= 3505;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S3522;
      end
      test_b1_S3522: begin
        IMAGE_addr <= 3506;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3512;
        test_state <= test_b1_S3523;
      end
      test_b1_S3523: begin
        IMAGE_addr <= 3507;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S3524;
      end
      test_b1_S3524: begin
        IMAGE_addr <= 3508;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S3525;
      end
      test_b1_S3525: begin
        IMAGE_addr <= 3509;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 107;
        test_state <= test_b1_S3526;
      end
      test_b1_S3526: begin
        IMAGE_addr <= 3510;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S3527;
      end
      test_b1_S3527: begin
        IMAGE_addr <= 3511;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3528;
      end
      test_b1_S3528: begin
        IMAGE_addr <= 3512;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3529;
      end
      test_b1_S3529: begin
        IMAGE_addr <= 3513;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3530;
      end
      test_b1_S3530: begin
        IMAGE_addr <= 3514;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S3531;
      end
      test_b1_S3531: begin
        IMAGE_addr <= 3515;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S3532;
      end
      test_b1_S3532: begin
        IMAGE_addr <= 3516;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3526;
        test_state <= test_b1_S3533;
      end
      test_b1_S3533: begin
        IMAGE_addr <= 3517;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S3534;
      end
      test_b1_S3534: begin
        IMAGE_addr <= 3518;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3523;
        test_state <= test_b1_S3535;
      end
      test_b1_S3535: begin
        IMAGE_addr <= 3519;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S3536;
      end
      test_b1_S3536: begin
        IMAGE_addr <= 3520;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 691;
        test_state <= test_b1_S3537;
      end
      test_b1_S3537: begin
        IMAGE_addr <= 3521;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 306;
        test_state <= test_b1_S3538;
      end
      test_b1_S3538: begin
        IMAGE_addr <= 3522;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3539;
      end
      test_b1_S3539: begin
        IMAGE_addr <= 3523;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 766;
        test_state <= test_b1_S3540;
      end
      test_b1_S3540: begin
        IMAGE_addr <= 3524;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 213;
        test_state <= test_b1_S3541;
      end
      test_b1_S3541: begin
        IMAGE_addr <= 3525;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3542;
      end
      test_b1_S3542: begin
        IMAGE_addr <= 3526;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 766;
        test_state <= test_b1_S3543;
      end
      test_b1_S3543: begin
        IMAGE_addr <= 3527;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 310;
        test_state <= test_b1_S3544;
      end
      test_b1_S3544: begin
        IMAGE_addr <= 3528;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S3545;
      end
      test_b1_S3545: begin
        IMAGE_addr <= 3529;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 708;
        test_state <= test_b1_S3546;
      end
      test_b1_S3546: begin
        IMAGE_addr <= 3530;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 306;
        test_state <= test_b1_S3547;
      end
      test_b1_S3547: begin
        IMAGE_addr <= 3531;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3548;
      end
      test_b1_S3548: begin
        IMAGE_addr <= 3532;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3549;
      end
      test_b1_S3549: begin
        IMAGE_addr <= 3533;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3504;
        test_state <= test_b1_S3550;
      end
      test_b1_S3550: begin
        IMAGE_addr <= 3534;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S3551;
      end
      test_b1_S3551: begin
        IMAGE_addr <= 3535;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3539;
        test_state <= test_b1_S3552;
      end
      test_b1_S3552: begin
        IMAGE_addr <= 3536;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 98;
        test_state <= test_b1_S3553;
      end
      test_b1_S3553: begin
        IMAGE_addr <= 3537;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S3554;
      end
      test_b1_S3554: begin
        IMAGE_addr <= 3538;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3555;
      end
      test_b1_S3555: begin
        IMAGE_addr <= 3539;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3556;
      end
      test_b1_S3556: begin
        IMAGE_addr <= 3540;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3557;
      end
      test_b1_S3557: begin
        IMAGE_addr <= 3541;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S3558;
      end
      test_b1_S3558: begin
        IMAGE_addr <= 3542;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 774;
        test_state <= test_b1_S3559;
      end
      test_b1_S3559: begin
        IMAGE_addr <= 3543;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 766;
        test_state <= test_b1_S3560;
      end
      test_b1_S3560: begin
        IMAGE_addr <= 3544;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 183;
        test_state <= test_b1_S3561;
      end
      test_b1_S3561: begin
        IMAGE_addr <= 3545;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3562;
      end
      test_b1_S3562: begin
        IMAGE_addr <= 3546;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3563;
      end
      test_b1_S3563: begin
        IMAGE_addr <= 3547;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3533;
        test_state <= test_b1_S3564;
      end
      test_b1_S3564: begin
        IMAGE_addr <= 3548;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S3565;
      end
      test_b1_S3565: begin
        IMAGE_addr <= 3549;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3554;
        test_state <= test_b1_S3566;
      end
      test_b1_S3566: begin
        IMAGE_addr <= 3550;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 98;
        test_state <= test_b1_S3567;
      end
      test_b1_S3567: begin
        IMAGE_addr <= 3551;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S3568;
      end
      test_b1_S3568: begin
        IMAGE_addr <= 3552;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 42;
        test_state <= test_b1_S3569;
      end
      test_b1_S3569: begin
        IMAGE_addr <= 3553;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3570;
      end
      test_b1_S3570: begin
        IMAGE_addr <= 3554;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3571;
      end
      test_b1_S3571: begin
        IMAGE_addr <= 3555;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3572;
      end
      test_b1_S3572: begin
        IMAGE_addr <= 3556;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S3573;
      end
      test_b1_S3573: begin
        IMAGE_addr <= 3557;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 766;
        test_state <= test_b1_S3574;
      end
      test_b1_S3574: begin
        IMAGE_addr <= 3558;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 766;
        test_state <= test_b1_S3575;
      end
      test_b1_S3575: begin
        IMAGE_addr <= 3559;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 183;
        test_state <= test_b1_S3576;
      end
      test_b1_S3576: begin
        IMAGE_addr <= 3560;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3577;
      end
      test_b1_S3577: begin
        IMAGE_addr <= 3561;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3578;
      end
      test_b1_S3578: begin
        IMAGE_addr <= 3562;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3547;
        test_state <= test_b1_S3579;
      end
      test_b1_S3579: begin
        IMAGE_addr <= 3563;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S3580;
      end
      test_b1_S3580: begin
        IMAGE_addr <= 3564;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3569;
        test_state <= test_b1_S3581;
      end
      test_b1_S3581: begin
        IMAGE_addr <= 3565;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 98;
        test_state <= test_b1_S3582;
      end
      test_b1_S3582: begin
        IMAGE_addr <= 3566;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S3583;
      end
      test_b1_S3583: begin
        IMAGE_addr <= 3567;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 64;
        test_state <= test_b1_S3584;
      end
      test_b1_S3584: begin
        IMAGE_addr <= 3568;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3585;
      end
      test_b1_S3585: begin
        IMAGE_addr <= 3569;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3586;
      end
      test_b1_S3586: begin
        IMAGE_addr <= 3570;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3587;
      end
      test_b1_S3587: begin
        IMAGE_addr <= 3571;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S3588;
      end
      test_b1_S3588: begin
        IMAGE_addr <= 3572;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3554;
        test_state <= test_b1_S3589;
      end
      test_b1_S3589: begin
        IMAGE_addr <= 3573;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3590;
      end
      test_b1_S3590: begin
        IMAGE_addr <= 3574;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3591;
      end
      test_b1_S3591: begin
        IMAGE_addr <= 3575;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3562;
        test_state <= test_b1_S3592;
      end
      test_b1_S3592: begin
        IMAGE_addr <= 3576;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S3593;
      end
      test_b1_S3593: begin
        IMAGE_addr <= 3577;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3582;
        test_state <= test_b1_S3594;
      end
      test_b1_S3594: begin
        IMAGE_addr <= 3578;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S3595;
      end
      test_b1_S3595: begin
        IMAGE_addr <= 3579;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S3596;
      end
      test_b1_S3596: begin
        IMAGE_addr <= 3580;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S3597;
      end
      test_b1_S3597: begin
        IMAGE_addr <= 3581;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3598;
      end
      test_b1_S3598: begin
        IMAGE_addr <= 3582;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3599;
      end
      test_b1_S3599: begin
        IMAGE_addr <= 3583;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3600;
      end
      test_b1_S3600: begin
        IMAGE_addr <= 3584;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S3601;
      end
      test_b1_S3601: begin
        IMAGE_addr <= 3585;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3591;
        test_state <= test_b1_S3602;
      end
      test_b1_S3602: begin
        IMAGE_addr <= 3586;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S3603;
      end
      test_b1_S3603: begin
        IMAGE_addr <= 3587;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 774;
        test_state <= test_b1_S3604;
      end
      test_b1_S3604: begin
        IMAGE_addr <= 3588;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 766;
        test_state <= test_b1_S3605;
      end
      test_b1_S3605: begin
        IMAGE_addr <= 3589;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 774;
        test_state <= test_b1_S3606;
      end
      test_b1_S3606: begin
        IMAGE_addr <= 3590;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3607;
      end
      test_b1_S3607: begin
        IMAGE_addr <= 3591;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 766;
        test_state <= test_b1_S3608;
      end
      test_b1_S3608: begin
        IMAGE_addr <= 3592;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 183;
        test_state <= test_b1_S3609;
      end
      test_b1_S3609: begin
        IMAGE_addr <= 3593;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3610;
      end
      test_b1_S3610: begin
        IMAGE_addr <= 3594;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3611;
      end
      test_b1_S3611: begin
        IMAGE_addr <= 3595;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3575;
        test_state <= test_b1_S3612;
      end
      test_b1_S3612: begin
        IMAGE_addr <= 3596;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S3613;
      end
      test_b1_S3613: begin
        IMAGE_addr <= 3597;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3603;
        test_state <= test_b1_S3614;
      end
      test_b1_S3614: begin
        IMAGE_addr <= 3598;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S3615;
      end
      test_b1_S3615: begin
        IMAGE_addr <= 3599;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S3616;
      end
      test_b1_S3616: begin
        IMAGE_addr <= 3600;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S3617;
      end
      test_b1_S3617: begin
        IMAGE_addr <= 3601;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 42;
        test_state <= test_b1_S3618;
      end
      test_b1_S3618: begin
        IMAGE_addr <= 3602;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3619;
      end
      test_b1_S3619: begin
        IMAGE_addr <= 3603;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3620;
      end
      test_b1_S3620: begin
        IMAGE_addr <= 3604;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3621;
      end
      test_b1_S3621: begin
        IMAGE_addr <= 3605;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S3622;
      end
      test_b1_S3622: begin
        IMAGE_addr <= 3606;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3617;
        test_state <= test_b1_S3623;
      end
      test_b1_S3623: begin
        IMAGE_addr <= 3607;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S3624;
      end
      test_b1_S3624: begin
        IMAGE_addr <= 3608;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3614;
        test_state <= test_b1_S3625;
      end
      test_b1_S3625: begin
        IMAGE_addr <= 3609;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S3626;
      end
      test_b1_S3626: begin
        IMAGE_addr <= 3610;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S3627;
      end
      test_b1_S3627: begin
        IMAGE_addr <= 3611;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 766;
        test_state <= test_b1_S3628;
      end
      test_b1_S3628: begin
        IMAGE_addr <= 3612;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 766;
        test_state <= test_b1_S3629;
      end
      test_b1_S3629: begin
        IMAGE_addr <= 3613;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3630;
      end
      test_b1_S3630: begin
        IMAGE_addr <= 3614;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 766;
        test_state <= test_b1_S3631;
      end
      test_b1_S3631: begin
        IMAGE_addr <= 3615;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 766;
        test_state <= test_b1_S3632;
      end
      test_b1_S3632: begin
        IMAGE_addr <= 3616;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3633;
      end
      test_b1_S3633: begin
        IMAGE_addr <= 3617;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 766;
        test_state <= test_b1_S3634;
      end
      test_b1_S3634: begin
        IMAGE_addr <= 3618;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 183;
        test_state <= test_b1_S3635;
      end
      test_b1_S3635: begin
        IMAGE_addr <= 3619;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3636;
      end
      test_b1_S3636: begin
        IMAGE_addr <= 3620;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3637;
      end
      test_b1_S3637: begin
        IMAGE_addr <= 3621;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3595;
        test_state <= test_b1_S3638;
      end
      test_b1_S3638: begin
        IMAGE_addr <= 3622;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S3639;
      end
      test_b1_S3639: begin
        IMAGE_addr <= 3623;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3629;
        test_state <= test_b1_S3640;
      end
      test_b1_S3640: begin
        IMAGE_addr <= 3624;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S3641;
      end
      test_b1_S3641: begin
        IMAGE_addr <= 3625;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S3642;
      end
      test_b1_S3642: begin
        IMAGE_addr <= 3626;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S3643;
      end
      test_b1_S3643: begin
        IMAGE_addr <= 3627;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 64;
        test_state <= test_b1_S3644;
      end
      test_b1_S3644: begin
        IMAGE_addr <= 3628;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3645;
      end
      test_b1_S3645: begin
        IMAGE_addr <= 3629;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3646;
      end
      test_b1_S3646: begin
        IMAGE_addr <= 3630;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3647;
      end
      test_b1_S3647: begin
        IMAGE_addr <= 3631;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S3648;
      end
      test_b1_S3648: begin
        IMAGE_addr <= 3632;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S3649;
      end
      test_b1_S3649: begin
        IMAGE_addr <= 3633;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3603;
        test_state <= test_b1_S3650;
      end
      test_b1_S3650: begin
        IMAGE_addr <= 3634;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3651;
      end
      test_b1_S3651: begin
        IMAGE_addr <= 3635;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3652;
      end
      test_b1_S3652: begin
        IMAGE_addr <= 3636;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3621;
        test_state <= test_b1_S3653;
      end
      test_b1_S3653: begin
        IMAGE_addr <= 3637;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S3654;
      end
      test_b1_S3654: begin
        IMAGE_addr <= 3638;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3644;
        test_state <= test_b1_S3655;
      end
      test_b1_S3655: begin
        IMAGE_addr <= 3639;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 99;
        test_state <= test_b1_S3656;
      end
      test_b1_S3656: begin
        IMAGE_addr <= 3640;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 111;
        test_state <= test_b1_S3657;
      end
      test_b1_S3657: begin
        IMAGE_addr <= 3641;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 110;
        test_state <= test_b1_S3658;
      end
      test_b1_S3658: begin
        IMAGE_addr <= 3642;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S3659;
      end
      test_b1_S3659: begin
        IMAGE_addr <= 3643;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3660;
      end
      test_b1_S3660: begin
        IMAGE_addr <= 3644;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3661;
      end
      test_b1_S3661: begin
        IMAGE_addr <= 3645;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3662;
      end
      test_b1_S3662: begin
        IMAGE_addr <= 3646;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5;
        test_state <= test_b1_S3663;
      end
      test_b1_S3663: begin
        IMAGE_addr <= 3647;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5;
        test_state <= test_b1_S3664;
      end
      test_b1_S3664: begin
        IMAGE_addr <= 3648;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S3665;
      end
      test_b1_S3665: begin
        IMAGE_addr <= 3649;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 691;
        test_state <= test_b1_S3666;
      end
      test_b1_S3666: begin
        IMAGE_addr <= 3650;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 306;
        test_state <= test_b1_S3667;
      end
      test_b1_S3667: begin
        IMAGE_addr <= 3651;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6;
        test_state <= test_b1_S3668;
      end
      test_b1_S3668: begin
        IMAGE_addr <= 3652;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6;
        test_state <= test_b1_S3669;
      end
      test_b1_S3669: begin
        IMAGE_addr <= 3653;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S3670;
      end
      test_b1_S3670: begin
        IMAGE_addr <= 3654;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 310;
        test_state <= test_b1_S3671;
      end
      test_b1_S3671: begin
        IMAGE_addr <= 3655;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3569;
        test_state <= test_b1_S3672;
      end
      test_b1_S3672: begin
        IMAGE_addr <= 3656;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S3673;
      end
      test_b1_S3673: begin
        IMAGE_addr <= 3657;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 708;
        test_state <= test_b1_S3674;
      end
      test_b1_S3674: begin
        IMAGE_addr <= 3658;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 306;
        test_state <= test_b1_S3675;
      end
      test_b1_S3675: begin
        IMAGE_addr <= 3659;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3676;
      end
      test_b1_S3676: begin
        IMAGE_addr <= 3660;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3677;
      end
      test_b1_S3677: begin
        IMAGE_addr <= 3661;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3636;
        test_state <= test_b1_S3678;
      end
      test_b1_S3678: begin
        IMAGE_addr <= 3662;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S3679;
      end
      test_b1_S3679: begin
        IMAGE_addr <= 3663;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3673;
        test_state <= test_b1_S3680;
      end
      test_b1_S3680: begin
        IMAGE_addr <= 3664;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 112;
        test_state <= test_b1_S3681;
      end
      test_b1_S3681: begin
        IMAGE_addr <= 3665;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S3682;
      end
      test_b1_S3682: begin
        IMAGE_addr <= 3666;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S3683;
      end
      test_b1_S3683: begin
        IMAGE_addr <= 3667;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S3684;
      end
      test_b1_S3684: begin
        IMAGE_addr <= 3668;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S3685;
      end
      test_b1_S3685: begin
        IMAGE_addr <= 3669;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S3686;
      end
      test_b1_S3686: begin
        IMAGE_addr <= 3670;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 118;
        test_state <= test_b1_S3687;
      end
      test_b1_S3687: begin
        IMAGE_addr <= 3671;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S3688;
      end
      test_b1_S3688: begin
        IMAGE_addr <= 3672;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3689;
      end
      test_b1_S3689: begin
        IMAGE_addr <= 3673;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3690;
      end
      test_b1_S3690: begin
        IMAGE_addr <= 3674;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3691;
      end
      test_b1_S3691: begin
        IMAGE_addr <= 3675;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S3692;
      end
      test_b1_S3692: begin
        IMAGE_addr <= 3676;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S3693;
      end
      test_b1_S3693: begin
        IMAGE_addr <= 3677;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 72;
        test_state <= test_b1_S3694;
      end
      test_b1_S3694: begin
        IMAGE_addr <= 3678;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 774;
        test_state <= test_b1_S3695;
      end
      test_b1_S3695: begin
        IMAGE_addr <= 3679;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S3696;
      end
      test_b1_S3696: begin
        IMAGE_addr <= 3680;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3685;
        test_state <= test_b1_S3697;
      end
      test_b1_S3697: begin
        IMAGE_addr <= 3681;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S3698;
      end
      test_b1_S3698: begin
        IMAGE_addr <= 3682;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 183;
        test_state <= test_b1_S3699;
      end
      test_b1_S3699: begin
        IMAGE_addr <= 3683;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 766;
        test_state <= test_b1_S3700;
      end
      test_b1_S3700: begin
        IMAGE_addr <= 3684;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3701;
      end
      test_b1_S3701: begin
        IMAGE_addr <= 3685;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 766;
        test_state <= test_b1_S3702;
      end
      test_b1_S3702: begin
        IMAGE_addr <= 3686;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S3703;
      end
      test_b1_S3703: begin
        IMAGE_addr <= 3687;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3704;
      end
      test_b1_S3704: begin
        IMAGE_addr <= 3688;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3705;
      end
      test_b1_S3705: begin
        IMAGE_addr <= 3689;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3661;
        test_state <= test_b1_S3706;
      end
      test_b1_S3706: begin
        IMAGE_addr <= 3690;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S3707;
      end
      test_b1_S3707: begin
        IMAGE_addr <= 3691;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3697;
        test_state <= test_b1_S3708;
      end
      test_b1_S3708: begin
        IMAGE_addr <= 3692;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 119;
        test_state <= test_b1_S3709;
      end
      test_b1_S3709: begin
        IMAGE_addr <= 3693;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 104;
        test_state <= test_b1_S3710;
      end
      test_b1_S3710: begin
        IMAGE_addr <= 3694;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S3711;
      end
      test_b1_S3711: begin
        IMAGE_addr <= 3695;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 110;
        test_state <= test_b1_S3712;
      end
      test_b1_S3712: begin
        IMAGE_addr <= 3696;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3713;
      end
      test_b1_S3713: begin
        IMAGE_addr <= 3697;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3714;
      end
      test_b1_S3714: begin
        IMAGE_addr <= 3698;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3715;
      end
      test_b1_S3715: begin
        IMAGE_addr <= 3699;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S3716;
      end
      test_b1_S3716: begin
        IMAGE_addr <= 3700;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3705;
        test_state <= test_b1_S3717;
      end
      test_b1_S3717: begin
        IMAGE_addr <= 3701;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 132;
        test_state <= test_b1_S3718;
      end
      test_b1_S3718: begin
        IMAGE_addr <= 3702;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S3719;
      end
      test_b1_S3719: begin
        IMAGE_addr <= 3703;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 183;
        test_state <= test_b1_S3720;
      end
      test_b1_S3720: begin
        IMAGE_addr <= 3704;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3721;
      end
      test_b1_S3721: begin
        IMAGE_addr <= 3705;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 766;
        test_state <= test_b1_S3722;
      end
      test_b1_S3722: begin
        IMAGE_addr <= 3706;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S3723;
      end
      test_b1_S3723: begin
        IMAGE_addr <= 3707;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S3724;
      end
      test_b1_S3724: begin
        IMAGE_addr <= 3708;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3713;
        test_state <= test_b1_S3725;
      end
      test_b1_S3725: begin
        IMAGE_addr <= 3709;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 183;
        test_state <= test_b1_S3726;
      end
      test_b1_S3726: begin
        IMAGE_addr <= 3710;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S3727;
      end
      test_b1_S3727: begin
        IMAGE_addr <= 3711;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4294967295;
        test_state <= test_b1_S3728;
      end
      test_b1_S3728: begin
        IMAGE_addr <= 3712;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3729;
      end
      test_b1_S3729: begin
        IMAGE_addr <= 3713;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S3730;
      end
      test_b1_S3730: begin
        IMAGE_addr <= 3714;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3719;
        test_state <= test_b1_S3731;
      end
      test_b1_S3731: begin
        IMAGE_addr <= 3715;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S3732;
      end
      test_b1_S3732: begin
        IMAGE_addr <= 3716;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S3733;
      end
      test_b1_S3733: begin
        IMAGE_addr <= 3717;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3734;
      end
      test_b1_S3734: begin
        IMAGE_addr <= 3718;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3735;
      end
      test_b1_S3735: begin
        IMAGE_addr <= 3719;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 732;
        test_state <= test_b1_S3736;
      end
      test_b1_S3736: begin
        IMAGE_addr <= 3720;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 25;
        test_state <= test_b1_S3737;
      end
      test_b1_S3737: begin
        IMAGE_addr <= 3721;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6;
        test_state <= test_b1_S3738;
      end
      test_b1_S3738: begin
        IMAGE_addr <= 3722;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S3739;
      end
      test_b1_S3739: begin
        IMAGE_addr <= 3723;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S3740;
      end
      test_b1_S3740: begin
        IMAGE_addr <= 3724;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3741;
      end
      test_b1_S3741: begin
        IMAGE_addr <= 3725;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3742;
      end
      test_b1_S3742: begin
        IMAGE_addr <= 3726;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3689;
        test_state <= test_b1_S3743;
      end
      test_b1_S3743: begin
        IMAGE_addr <= 3727;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S3744;
      end
      test_b1_S3744: begin
        IMAGE_addr <= 3728;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3735;
        test_state <= test_b1_S3745;
      end
      test_b1_S3745: begin
        IMAGE_addr <= 3729;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 119;
        test_state <= test_b1_S3746;
      end
      test_b1_S3746: begin
        IMAGE_addr <= 3730;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 104;
        test_state <= test_b1_S3747;
      end
      test_b1_S3747: begin
        IMAGE_addr <= 3731;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S3748;
      end
      test_b1_S3748: begin
        IMAGE_addr <= 3732;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 110;
        test_state <= test_b1_S3749;
      end
      test_b1_S3749: begin
        IMAGE_addr <= 3733;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 100;
        test_state <= test_b1_S3750;
      end
      test_b1_S3750: begin
        IMAGE_addr <= 3734;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3751;
      end
      test_b1_S3751: begin
        IMAGE_addr <= 3735;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3752;
      end
      test_b1_S3752: begin
        IMAGE_addr <= 3736;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3753;
      end
      test_b1_S3753: begin
        IMAGE_addr <= 3737;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S3754;
      end
      test_b1_S3754: begin
        IMAGE_addr <= 3738;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3743;
        test_state <= test_b1_S3755;
      end
      test_b1_S3755: begin
        IMAGE_addr <= 3739;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 132;
        test_state <= test_b1_S3756;
      end
      test_b1_S3756: begin
        IMAGE_addr <= 3740;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S3757;
      end
      test_b1_S3757: begin
        IMAGE_addr <= 3741;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 183;
        test_state <= test_b1_S3758;
      end
      test_b1_S3758: begin
        IMAGE_addr <= 3742;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3759;
      end
      test_b1_S3759: begin
        IMAGE_addr <= 3743;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 766;
        test_state <= test_b1_S3760;
      end
      test_b1_S3760: begin
        IMAGE_addr <= 3744;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S3761;
      end
      test_b1_S3761: begin
        IMAGE_addr <= 3745;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S3762;
      end
      test_b1_S3762: begin
        IMAGE_addr <= 3746;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3752;
        test_state <= test_b1_S3763;
      end
      test_b1_S3763: begin
        IMAGE_addr <= 3747;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2577;
        test_state <= test_b1_S3764;
      end
      test_b1_S3764: begin
        IMAGE_addr <= 3748;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 183;
        test_state <= test_b1_S3765;
      end
      test_b1_S3765: begin
        IMAGE_addr <= 3749;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S3766;
      end
      test_b1_S3766: begin
        IMAGE_addr <= 3750;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4294967295;
        test_state <= test_b1_S3767;
      end
      test_b1_S3767: begin
        IMAGE_addr <= 3751;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3768;
      end
      test_b1_S3768: begin
        IMAGE_addr <= 3752;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S3769;
      end
      test_b1_S3769: begin
        IMAGE_addr <= 3753;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3758;
        test_state <= test_b1_S3770;
      end
      test_b1_S3770: begin
        IMAGE_addr <= 3754;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S3771;
      end
      test_b1_S3771: begin
        IMAGE_addr <= 3755;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S3772;
      end
      test_b1_S3772: begin
        IMAGE_addr <= 3756;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3773;
      end
      test_b1_S3773: begin
        IMAGE_addr <= 3757;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3774;
      end
      test_b1_S3774: begin
        IMAGE_addr <= 3758;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 732;
        test_state <= test_b1_S3775;
      end
      test_b1_S3775: begin
        IMAGE_addr <= 3759;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 25;
        test_state <= test_b1_S3776;
      end
      test_b1_S3776: begin
        IMAGE_addr <= 3760;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6;
        test_state <= test_b1_S3777;
      end
      test_b1_S3777: begin
        IMAGE_addr <= 3761;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S3778;
      end
      test_b1_S3778: begin
        IMAGE_addr <= 3762;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S3779;
      end
      test_b1_S3779: begin
        IMAGE_addr <= 3763;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3780;
      end
      test_b1_S3780: begin
        IMAGE_addr <= 3764;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3781;
      end
      test_b1_S3781: begin
        IMAGE_addr <= 3765;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3726;
        test_state <= test_b1_S3782;
      end
      test_b1_S3782: begin
        IMAGE_addr <= 3766;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3283;
        test_state <= test_b1_S3783;
      end
      test_b1_S3783: begin
        IMAGE_addr <= 3767;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3772;
        test_state <= test_b1_S3784;
      end
      test_b1_S3784: begin
        IMAGE_addr <= 3768;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 102;
        test_state <= test_b1_S3785;
      end
      test_b1_S3785: begin
        IMAGE_addr <= 3769;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 111;
        test_state <= test_b1_S3786;
      end
      test_b1_S3786: begin
        IMAGE_addr <= 3770;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S3787;
      end
      test_b1_S3787: begin
        IMAGE_addr <= 3771;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3788;
      end
      test_b1_S3788: begin
        IMAGE_addr <= 3772;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 206;
        test_state <= test_b1_S3789;
      end
      test_b1_S3789: begin
        IMAGE_addr <= 3773;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S3790;
      end
      test_b1_S3790: begin
        IMAGE_addr <= 3774;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 252;
        test_state <= test_b1_S3791;
      end
      test_b1_S3791: begin
        IMAGE_addr <= 3775;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3283;
        test_state <= test_b1_S3792;
      end
      test_b1_S3792: begin
        IMAGE_addr <= 3776;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3793;
      end
      test_b1_S3793: begin
        IMAGE_addr <= 3777;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3794;
      end
      test_b1_S3794: begin
        IMAGE_addr <= 3778;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3765;
        test_state <= test_b1_S3795;
      end
      test_b1_S3795: begin
        IMAGE_addr <= 3779;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3283;
        test_state <= test_b1_S3796;
      end
      test_b1_S3796: begin
        IMAGE_addr <= 3780;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3786;
        test_state <= test_b1_S3797;
      end
      test_b1_S3797: begin
        IMAGE_addr <= 3781;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 110;
        test_state <= test_b1_S3798;
      end
      test_b1_S3798: begin
        IMAGE_addr <= 3782;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S3799;
      end
      test_b1_S3799: begin
        IMAGE_addr <= 3783;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 120;
        test_state <= test_b1_S3800;
      end
      test_b1_S3800: begin
        IMAGE_addr <= 3784;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S3801;
      end
      test_b1_S3801: begin
        IMAGE_addr <= 3785;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3802;
      end
      test_b1_S3802: begin
        IMAGE_addr <= 3786;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S3803;
      end
      test_b1_S3803: begin
        IMAGE_addr <= 3787;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 259;
        test_state <= test_b1_S3804;
      end
      test_b1_S3804: begin
        IMAGE_addr <= 3788;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3283;
        test_state <= test_b1_S3805;
      end
      test_b1_S3805: begin
        IMAGE_addr <= 3789;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S3806;
      end
      test_b1_S3806: begin
        IMAGE_addr <= 3790;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7;
        test_state <= test_b1_S3807;
      end
      test_b1_S3807: begin
        IMAGE_addr <= 3791;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 213;
        test_state <= test_b1_S3808;
      end
      test_b1_S3808: begin
        IMAGE_addr <= 3792;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 213;
        test_state <= test_b1_S3809;
      end
      test_b1_S3809: begin
        IMAGE_addr <= 3793;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3810;
      end
      test_b1_S3810: begin
        IMAGE_addr <= 3794;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3811;
      end
      test_b1_S3811: begin
        IMAGE_addr <= 3795;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3778;
        test_state <= test_b1_S3812;
      end
      test_b1_S3812: begin
        IMAGE_addr <= 3796;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S3813;
      end
      test_b1_S3813: begin
        IMAGE_addr <= 3797;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3800;
        test_state <= test_b1_S3814;
      end
      test_b1_S3814: begin
        IMAGE_addr <= 3798;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S3815;
      end
      test_b1_S3815: begin
        IMAGE_addr <= 3799;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3816;
      end
      test_b1_S3816: begin
        IMAGE_addr <= 3800;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6;
        test_state <= test_b1_S3817;
      end
      test_b1_S3817: begin
        IMAGE_addr <= 3801;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6;
        test_state <= test_b1_S3818;
      end
      test_b1_S3818: begin
        IMAGE_addr <= 3802;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6;
        test_state <= test_b1_S3819;
      end
      test_b1_S3819: begin
        IMAGE_addr <= 3803;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 132;
        test_state <= test_b1_S3820;
      end
      test_b1_S3820: begin
        IMAGE_addr <= 3804;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 132;
        test_state <= test_b1_S3821;
      end
      test_b1_S3821: begin
        IMAGE_addr <= 3805;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5;
        test_state <= test_b1_S3822;
      end
      test_b1_S3822: begin
        IMAGE_addr <= 3806;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5;
        test_state <= test_b1_S3823;
      end
      test_b1_S3823: begin
        IMAGE_addr <= 3807;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S3824;
      end
      test_b1_S3824: begin
        IMAGE_addr <= 3808;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 17;
        test_state <= test_b1_S3825;
      end
      test_b1_S3825: begin
        IMAGE_addr <= 3809;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S3826;
      end
      test_b1_S3826: begin
        IMAGE_addr <= 3810;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5;
        test_state <= test_b1_S3827;
      end
      test_b1_S3827: begin
        IMAGE_addr <= 3811;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3828;
      end
      test_b1_S3828: begin
        IMAGE_addr <= 3812;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3829;
      end
      test_b1_S3829: begin
        IMAGE_addr <= 3813;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3795;
        test_state <= test_b1_S3830;
      end
      test_b1_S3830: begin
        IMAGE_addr <= 3814;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3283;
        test_state <= test_b1_S3831;
      end
      test_b1_S3831: begin
        IMAGE_addr <= 3815;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3821;
        test_state <= test_b1_S3832;
      end
      test_b1_S3832: begin
        IMAGE_addr <= 3816;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S3833;
      end
      test_b1_S3833: begin
        IMAGE_addr <= 3817;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 111;
        test_state <= test_b1_S3834;
      end
      test_b1_S3834: begin
        IMAGE_addr <= 3818;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S3835;
      end
      test_b1_S3835: begin
        IMAGE_addr <= 3819;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S3836;
      end
      test_b1_S3836: begin
        IMAGE_addr <= 3820;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3837;
      end
      test_b1_S3837: begin
        IMAGE_addr <= 3821;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S3838;
      end
      test_b1_S3838: begin
        IMAGE_addr <= 3822;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 259;
        test_state <= test_b1_S3839;
      end
      test_b1_S3839: begin
        IMAGE_addr <= 3823;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3283;
        test_state <= test_b1_S3840;
      end
      test_b1_S3840: begin
        IMAGE_addr <= 3824;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S3841;
      end
      test_b1_S3841: begin
        IMAGE_addr <= 3825;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 32;
        test_state <= test_b1_S3842;
      end
      test_b1_S3842: begin
        IMAGE_addr <= 3826;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 323;
        test_state <= test_b1_S3843;
      end
      test_b1_S3843: begin
        IMAGE_addr <= 3827;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S3844;
      end
      test_b1_S3844: begin
        IMAGE_addr <= 3828;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 252;
        test_state <= test_b1_S3845;
      end
      test_b1_S3845: begin
        IMAGE_addr <= 3829;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3283;
        test_state <= test_b1_S3846;
      end
      test_b1_S3846: begin
        IMAGE_addr <= 3830;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3847;
      end
      test_b1_S3847: begin
        IMAGE_addr <= 3831;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3848;
      end
      test_b1_S3848: begin
        IMAGE_addr <= 3832;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3726;
        test_state <= test_b1_S3849;
      end
      test_b1_S3849: begin
        IMAGE_addr <= 3833;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S3850;
      end
      test_b1_S3850: begin
        IMAGE_addr <= 3834;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3841;
        test_state <= test_b1_S3851;
      end
      test_b1_S3851: begin
        IMAGE_addr <= 3835;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S3852;
      end
      test_b1_S3852: begin
        IMAGE_addr <= 3836;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S3853;
      end
      test_b1_S3853: begin
        IMAGE_addr <= 3837;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 109;
        test_state <= test_b1_S3854;
      end
      test_b1_S3854: begin
        IMAGE_addr <= 3838;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S3855;
      end
      test_b1_S3855: begin
        IMAGE_addr <= 3839;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S3856;
      end
      test_b1_S3856: begin
        IMAGE_addr <= 3840;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3857;
      end
      test_b1_S3857: begin
        IMAGE_addr <= 3841;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3858;
      end
      test_b1_S3858: begin
        IMAGE_addr <= 3842;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3859;
      end
      test_b1_S3859: begin
        IMAGE_addr <= 3843;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 132;
        test_state <= test_b1_S3860;
      end
      test_b1_S3860: begin
        IMAGE_addr <= 3844;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S3861;
      end
      test_b1_S3861: begin
        IMAGE_addr <= 3845;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S3862;
      end
      test_b1_S3862: begin
        IMAGE_addr <= 3846;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 806;
        test_state <= test_b1_S3863;
      end
      test_b1_S3863: begin
        IMAGE_addr <= 3847;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S3864;
      end
      test_b1_S3864: begin
        IMAGE_addr <= 3848;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3858;
        test_state <= test_b1_S3865;
      end
      test_b1_S3865: begin
        IMAGE_addr <= 3849;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S3866;
      end
      test_b1_S3866: begin
        IMAGE_addr <= 3850;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5;
        test_state <= test_b1_S3867;
      end
      test_b1_S3867: begin
        IMAGE_addr <= 3851;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S3868;
      end
      test_b1_S3868: begin
        IMAGE_addr <= 3852;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 766;
        test_state <= test_b1_S3869;
      end
      test_b1_S3869: begin
        IMAGE_addr <= 3853;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6;
        test_state <= test_b1_S3870;
      end
      test_b1_S3870: begin
        IMAGE_addr <= 3854;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7;
        test_state <= test_b1_S3871;
      end
      test_b1_S3871: begin
        IMAGE_addr <= 3855;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3850;
        test_state <= test_b1_S3872;
      end
      test_b1_S3872: begin
        IMAGE_addr <= 3856;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S3873;
      end
      test_b1_S3873: begin
        IMAGE_addr <= 3857;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3874;
      end
      test_b1_S3874: begin
        IMAGE_addr <= 3858;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S3875;
      end
      test_b1_S3875: begin
        IMAGE_addr <= 3859;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3863;
        test_state <= test_b1_S3876;
      end
      test_b1_S3876: begin
        IMAGE_addr <= 3860;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S3877;
      end
      test_b1_S3877: begin
        IMAGE_addr <= 3861;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S3878;
      end
      test_b1_S3878: begin
        IMAGE_addr <= 3862;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3879;
      end
      test_b1_S3879: begin
        IMAGE_addr <= 3863;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 732;
        test_state <= test_b1_S3880;
      end
      test_b1_S3880: begin
        IMAGE_addr <= 3864;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3881;
      end
      test_b1_S3881: begin
        IMAGE_addr <= 3865;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3882;
      end
      test_b1_S3882: begin
        IMAGE_addr <= 3866;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3832;
        test_state <= test_b1_S3883;
      end
      test_b1_S3883: begin
        IMAGE_addr <= 3867;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S3884;
      end
      test_b1_S3884: begin
        IMAGE_addr <= 3868;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3875;
        test_state <= test_b1_S3885;
      end
      test_b1_S3885: begin
        IMAGE_addr <= 3869;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S3886;
      end
      test_b1_S3886: begin
        IMAGE_addr <= 3870;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S3887;
      end
      test_b1_S3887: begin
        IMAGE_addr <= 3871;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S3888;
      end
      test_b1_S3888: begin
        IMAGE_addr <= 3872;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S3889;
      end
      test_b1_S3889: begin
        IMAGE_addr <= 3873;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 100;
        test_state <= test_b1_S3890;
      end
      test_b1_S3890: begin
        IMAGE_addr <= 3874;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3891;
      end
      test_b1_S3891: begin
        IMAGE_addr <= 3875;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3892;
      end
      test_b1_S3892: begin
        IMAGE_addr <= 3876;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3893;
      end
      test_b1_S3893: begin
        IMAGE_addr <= 3877;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 132;
        test_state <= test_b1_S3894;
      end
      test_b1_S3894: begin
        IMAGE_addr <= 3878;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S3895;
      end
      test_b1_S3895: begin
        IMAGE_addr <= 3879;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S3896;
      end
      test_b1_S3896: begin
        IMAGE_addr <= 3880;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 806;
        test_state <= test_b1_S3897;
      end
      test_b1_S3897: begin
        IMAGE_addr <= 3881;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S3898;
      end
      test_b1_S3898: begin
        IMAGE_addr <= 3882;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3896;
        test_state <= test_b1_S3899;
      end
      test_b1_S3899: begin
        IMAGE_addr <= 3883;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S3900;
      end
      test_b1_S3900: begin
        IMAGE_addr <= 3884;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5;
        test_state <= test_b1_S3901;
      end
      test_b1_S3901: begin
        IMAGE_addr <= 3885;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6;
        test_state <= test_b1_S3902;
      end
      test_b1_S3902: begin
        IMAGE_addr <= 3886;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S3903;
      end
      test_b1_S3903: begin
        IMAGE_addr <= 3887;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5;
        test_state <= test_b1_S3904;
      end
      test_b1_S3904: begin
        IMAGE_addr <= 3888;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S3905;
      end
      test_b1_S3905: begin
        IMAGE_addr <= 3889;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S3906;
      end
      test_b1_S3906: begin
        IMAGE_addr <= 3890;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 766;
        test_state <= test_b1_S3907;
      end
      test_b1_S3907: begin
        IMAGE_addr <= 3891;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6;
        test_state <= test_b1_S3908;
      end
      test_b1_S3908: begin
        IMAGE_addr <= 3892;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7;
        test_state <= test_b1_S3909;
      end
      test_b1_S3909: begin
        IMAGE_addr <= 3893;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3884;
        test_state <= test_b1_S3910;
      end
      test_b1_S3910: begin
        IMAGE_addr <= 3894;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S3911;
      end
      test_b1_S3911: begin
        IMAGE_addr <= 3895;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3912;
      end
      test_b1_S3912: begin
        IMAGE_addr <= 3896;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S3913;
      end
      test_b1_S3913: begin
        IMAGE_addr <= 3897;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3901;
        test_state <= test_b1_S3914;
      end
      test_b1_S3914: begin
        IMAGE_addr <= 3898;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S3915;
      end
      test_b1_S3915: begin
        IMAGE_addr <= 3899;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S3916;
      end
      test_b1_S3916: begin
        IMAGE_addr <= 3900;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3917;
      end
      test_b1_S3917: begin
        IMAGE_addr <= 3901;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 732;
        test_state <= test_b1_S3918;
      end
      test_b1_S3918: begin
        IMAGE_addr <= 3902;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3919;
      end
      test_b1_S3919: begin
        IMAGE_addr <= 3903;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3920;
      end
      test_b1_S3920: begin
        IMAGE_addr <= 3904;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3866;
        test_state <= test_b1_S3921;
      end
      test_b1_S3921: begin
        IMAGE_addr <= 3905;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S3922;
      end
      test_b1_S3922: begin
        IMAGE_addr <= 3906;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3912;
        test_state <= test_b1_S3923;
      end
      test_b1_S3923: begin
        IMAGE_addr <= 3907;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S3924;
      end
      test_b1_S3924: begin
        IMAGE_addr <= 3908;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S3925;
      end
      test_b1_S3925: begin
        IMAGE_addr <= 3909;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S3926;
      end
      test_b1_S3926: begin
        IMAGE_addr <= 3910;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S3927;
      end
      test_b1_S3927: begin
        IMAGE_addr <= 3911;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3928;
      end
      test_b1_S3928: begin
        IMAGE_addr <= 3912;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3929;
      end
      test_b1_S3929: begin
        IMAGE_addr <= 3913;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3930;
      end
      test_b1_S3930: begin
        IMAGE_addr <= 3914;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 132;
        test_state <= test_b1_S3931;
      end
      test_b1_S3931: begin
        IMAGE_addr <= 3915;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S3932;
      end
      test_b1_S3932: begin
        IMAGE_addr <= 3916;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S3933;
      end
      test_b1_S3933: begin
        IMAGE_addr <= 3917;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 806;
        test_state <= test_b1_S3934;
      end
      test_b1_S3934: begin
        IMAGE_addr <= 3918;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S3935;
      end
      test_b1_S3935: begin
        IMAGE_addr <= 3919;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3935;
        test_state <= test_b1_S3936;
      end
      test_b1_S3936: begin
        IMAGE_addr <= 3920;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S3937;
      end
      test_b1_S3937: begin
        IMAGE_addr <= 3921;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S3938;
      end
      test_b1_S3938: begin
        IMAGE_addr <= 3922;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5;
        test_state <= test_b1_S3939;
      end
      test_b1_S3939: begin
        IMAGE_addr <= 3923;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5;
        test_state <= test_b1_S3940;
      end
      test_b1_S3940: begin
        IMAGE_addr <= 3924;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3800;
        test_state <= test_b1_S3941;
      end
      test_b1_S3941: begin
        IMAGE_addr <= 3925;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S3942;
      end
      test_b1_S3942: begin
        IMAGE_addr <= 3926;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S3943;
      end
      test_b1_S3943: begin
        IMAGE_addr <= 3927;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 766;
        test_state <= test_b1_S3944;
      end
      test_b1_S3944: begin
        IMAGE_addr <= 3928;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6;
        test_state <= test_b1_S3945;
      end
      test_b1_S3945: begin
        IMAGE_addr <= 3929;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7;
        test_state <= test_b1_S3946;
      end
      test_b1_S3946: begin
        IMAGE_addr <= 3930;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3923;
        test_state <= test_b1_S3947;
      end
      test_b1_S3947: begin
        IMAGE_addr <= 3931;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6;
        test_state <= test_b1_S3948;
      end
      test_b1_S3948: begin
        IMAGE_addr <= 3932;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S3949;
      end
      test_b1_S3949: begin
        IMAGE_addr <= 3933;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S3950;
      end
      test_b1_S3950: begin
        IMAGE_addr <= 3934;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3951;
      end
      test_b1_S3951: begin
        IMAGE_addr <= 3935;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S3952;
      end
      test_b1_S3952: begin
        IMAGE_addr <= 3936;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3940;
        test_state <= test_b1_S3953;
      end
      test_b1_S3953: begin
        IMAGE_addr <= 3937;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S3954;
      end
      test_b1_S3954: begin
        IMAGE_addr <= 3938;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S3955;
      end
      test_b1_S3955: begin
        IMAGE_addr <= 3939;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3956;
      end
      test_b1_S3956: begin
        IMAGE_addr <= 3940;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 732;
        test_state <= test_b1_S3957;
      end
      test_b1_S3957: begin
        IMAGE_addr <= 3941;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3958;
      end
      test_b1_S3958: begin
        IMAGE_addr <= 3942;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3959;
      end
      test_b1_S3959: begin
        IMAGE_addr <= 3943;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3904;
        test_state <= test_b1_S3960;
      end
      test_b1_S3960: begin
        IMAGE_addr <= 3944;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S3961;
      end
      test_b1_S3961: begin
        IMAGE_addr <= 3945;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3951;
        test_state <= test_b1_S3962;
      end
      test_b1_S3962: begin
        IMAGE_addr <= 3946;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S3963;
      end
      test_b1_S3963: begin
        IMAGE_addr <= 3947;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S3964;
      end
      test_b1_S3964: begin
        IMAGE_addr <= 3948;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 99;
        test_state <= test_b1_S3965;
      end
      test_b1_S3965: begin
        IMAGE_addr <= 3949;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 104;
        test_state <= test_b1_S3966;
      end
      test_b1_S3966: begin
        IMAGE_addr <= 3950;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3967;
      end
      test_b1_S3967: begin
        IMAGE_addr <= 3951;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S3968;
      end
      test_b1_S3968: begin
        IMAGE_addr <= 3952;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3964;
        test_state <= test_b1_S3969;
      end
      test_b1_S3969: begin
        IMAGE_addr <= 3953;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S3970;
      end
      test_b1_S3970: begin
        IMAGE_addr <= 3954;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3961;
        test_state <= test_b1_S3971;
      end
      test_b1_S3971: begin
        IMAGE_addr <= 3955;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S3972;
      end
      test_b1_S3972: begin
        IMAGE_addr <= 3956;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S3973;
      end
      test_b1_S3973: begin
        IMAGE_addr <= 3957;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S3974;
      end
      test_b1_S3974: begin
        IMAGE_addr <= 3958;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 183;
        test_state <= test_b1_S3975;
      end
      test_b1_S3975: begin
        IMAGE_addr <= 3959;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 766;
        test_state <= test_b1_S3976;
      end
      test_b1_S3976: begin
        IMAGE_addr <= 3960;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3977;
      end
      test_b1_S3977: begin
        IMAGE_addr <= 3961;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 774;
        test_state <= test_b1_S3978;
      end
      test_b1_S3978: begin
        IMAGE_addr <= 3962;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 26;
        test_state <= test_b1_S3979;
      end
      test_b1_S3979: begin
        IMAGE_addr <= 3963;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3980;
      end
      test_b1_S3980: begin
        IMAGE_addr <= 3964;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3841;
        test_state <= test_b1_S3981;
      end
      test_b1_S3981: begin
        IMAGE_addr <= 3965;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S3982;
      end
      test_b1_S3982: begin
        IMAGE_addr <= 3966;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S3983;
      end
      test_b1_S3983: begin
        IMAGE_addr <= 3967;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3984;
      end
      test_b1_S3984: begin
        IMAGE_addr <= 3968;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S3985;
      end
      test_b1_S3985: begin
        IMAGE_addr <= 3969;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3943;
        test_state <= test_b1_S3986;
      end
      test_b1_S3986: begin
        IMAGE_addr <= 3970;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S3987;
      end
      test_b1_S3987: begin
        IMAGE_addr <= 3971;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3978;
        test_state <= test_b1_S3988;
      end
      test_b1_S3988: begin
        IMAGE_addr <= 3972;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S3989;
      end
      test_b1_S3989: begin
        IMAGE_addr <= 3973;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S3990;
      end
      test_b1_S3990: begin
        IMAGE_addr <= 3974;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S3991;
      end
      test_b1_S3991: begin
        IMAGE_addr <= 3975;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S3992;
      end
      test_b1_S3992: begin
        IMAGE_addr <= 3976;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 121;
        test_state <= test_b1_S3993;
      end
      test_b1_S3993: begin
        IMAGE_addr <= 3977;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S3994;
      end
      test_b1_S3994: begin
        IMAGE_addr <= 3978;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S3995;
      end
      test_b1_S3995: begin
        IMAGE_addr <= 3979;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 189;
        test_state <= test_b1_S3996;
      end
      test_b1_S3996: begin
        IMAGE_addr <= 3980;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S3997;
      end
      test_b1_S3997: begin
        IMAGE_addr <= 3981;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S3998;
      end
      test_b1_S3998: begin
        IMAGE_addr <= 3982;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S3999;
      end
      test_b1_S3999: begin
        IMAGE_addr <= 3983;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 830;
        test_state <= test_b1_S4000;
      end
      test_b1_S4000: begin
        IMAGE_addr <= 3984;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S4001;
      end
      test_b1_S4001: begin
        IMAGE_addr <= 3985;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3988;
        test_state <= test_b1_S4002;
      end
      test_b1_S4002: begin
        IMAGE_addr <= 3986;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3951;
        test_state <= test_b1_S4003;
      end
      test_b1_S4003: begin
        IMAGE_addr <= 3987;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4004;
      end
      test_b1_S4004: begin
        IMAGE_addr <= 3988;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S4005;
      end
      test_b1_S4005: begin
        IMAGE_addr <= 3989;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3993;
        test_state <= test_b1_S4006;
      end
      test_b1_S4006: begin
        IMAGE_addr <= 3990;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S4007;
      end
      test_b1_S4007: begin
        IMAGE_addr <= 3991;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S4008;
      end
      test_b1_S4008: begin
        IMAGE_addr <= 3992;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4009;
      end
      test_b1_S4009: begin
        IMAGE_addr <= 3993;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 732;
        test_state <= test_b1_S4010;
      end
      test_b1_S4010: begin
        IMAGE_addr <= 3994;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4011;
      end
      test_b1_S4011: begin
        IMAGE_addr <= 3995;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4012;
      end
      test_b1_S4012: begin
        IMAGE_addr <= 3996;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3969;
        test_state <= test_b1_S4013;
      end
      test_b1_S4013: begin
        IMAGE_addr <= 3997;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S4014;
      end
      test_b1_S4014: begin
        IMAGE_addr <= 3998;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4006;
        test_state <= test_b1_S4015;
      end
      test_b1_S4015: begin
        IMAGE_addr <= 3999;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 98;
        test_state <= test_b1_S4016;
      end
      test_b1_S4016: begin
        IMAGE_addr <= 4000;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 117;
        test_state <= test_b1_S4017;
      end
      test_b1_S4017: begin
        IMAGE_addr <= 4001;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 102;
        test_state <= test_b1_S4018;
      end
      test_b1_S4018: begin
        IMAGE_addr <= 4002;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 102;
        test_state <= test_b1_S4019;
      end
      test_b1_S4019: begin
        IMAGE_addr <= 4003;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S4020;
      end
      test_b1_S4020: begin
        IMAGE_addr <= 4004;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S4021;
      end
      test_b1_S4021: begin
        IMAGE_addr <= 4005;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4022;
      end
      test_b1_S4022: begin
        IMAGE_addr <= 4006;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2590;
        test_state <= test_b1_S4023;
      end
      test_b1_S4023: begin
        IMAGE_addr <= 4007;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2590;
        test_state <= test_b1_S4024;
      end
      test_b1_S4024: begin
        IMAGE_addr <= 4008;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3951;
        test_state <= test_b1_S4025;
      end
      test_b1_S4025: begin
        IMAGE_addr <= 4009;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4026;
      end
      test_b1_S4026: begin
        IMAGE_addr <= 4010;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4027;
      end
      test_b1_S4027: begin
        IMAGE_addr <= 4011;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3996;
        test_state <= test_b1_S4028;
      end
      test_b1_S4028: begin
        IMAGE_addr <= 4012;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S4029;
      end
      test_b1_S4029: begin
        IMAGE_addr <= 4013;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4019;
        test_state <= test_b1_S4030;
      end
      test_b1_S4030: begin
        IMAGE_addr <= 4014;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 108;
        test_state <= test_b1_S4031;
      end
      test_b1_S4031: begin
        IMAGE_addr <= 4015;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S4032;
      end
      test_b1_S4032: begin
        IMAGE_addr <= 4016;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S4033;
      end
      test_b1_S4033: begin
        IMAGE_addr <= 4017;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S4034;
      end
      test_b1_S4034: begin
        IMAGE_addr <= 4018;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4035;
      end
      test_b1_S4035: begin
        IMAGE_addr <= 4019;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S4036;
      end
      test_b1_S4036: begin
        IMAGE_addr <= 4020;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4036;
        test_state <= test_b1_S4037;
      end
      test_b1_S4037: begin
        IMAGE_addr <= 4021;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S4038;
      end
      test_b1_S4038: begin
        IMAGE_addr <= 4022;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 72;
        test_state <= test_b1_S4039;
      end
      test_b1_S4039: begin
        IMAGE_addr <= 4023;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 766;
        test_state <= test_b1_S4040;
      end
      test_b1_S4040: begin
        IMAGE_addr <= 4024;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 132;
        test_state <= test_b1_S4041;
      end
      test_b1_S4041: begin
        IMAGE_addr <= 4025;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 132;
        test_state <= test_b1_S4042;
      end
      test_b1_S4042: begin
        IMAGE_addr <= 4026;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S4043;
      end
      test_b1_S4043: begin
        IMAGE_addr <= 4027;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4032;
        test_state <= test_b1_S4044;
      end
      test_b1_S4044: begin
        IMAGE_addr <= 4028;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S4045;
      end
      test_b1_S4045: begin
        IMAGE_addr <= 4029;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 183;
        test_state <= test_b1_S4046;
      end
      test_b1_S4046: begin
        IMAGE_addr <= 4030;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 766;
        test_state <= test_b1_S4047;
      end
      test_b1_S4047: begin
        IMAGE_addr <= 4031;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4048;
      end
      test_b1_S4048: begin
        IMAGE_addr <= 4032;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 766;
        test_state <= test_b1_S4049;
      end
      test_b1_S4049: begin
        IMAGE_addr <= 4033;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 132;
        test_state <= test_b1_S4050;
      end
      test_b1_S4050: begin
        IMAGE_addr <= 4034;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S4051;
      end
      test_b1_S4051: begin
        IMAGE_addr <= 4035;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4052;
      end
      test_b1_S4052: begin
        IMAGE_addr <= 4036;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3433;
        test_state <= test_b1_S4053;
      end
      test_b1_S4053: begin
        IMAGE_addr <= 4037;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S4054;
      end
      test_b1_S4054: begin
        IMAGE_addr <= 4038;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S4055;
      end
      test_b1_S4055: begin
        IMAGE_addr <= 4039;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4056;
      end
      test_b1_S4056: begin
        IMAGE_addr <= 4040;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4057;
      end
      test_b1_S4057: begin
        IMAGE_addr <= 4041;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3904;
        test_state <= test_b1_S4058;
      end
      test_b1_S4058: begin
        IMAGE_addr <= 4042;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S4059;
      end
      test_b1_S4059: begin
        IMAGE_addr <= 4043;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4052;
        test_state <= test_b1_S4060;
      end
      test_b1_S4060: begin
        IMAGE_addr <= 4044;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 60;
        test_state <= test_b1_S4061;
      end
      test_b1_S4061: begin
        IMAGE_addr <= 4045;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S4062;
      end
      test_b1_S4062: begin
        IMAGE_addr <= 4046;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S4063;
      end
      test_b1_S4063: begin
        IMAGE_addr <= 4047;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 99;
        test_state <= test_b1_S4064;
      end
      test_b1_S4064: begin
        IMAGE_addr <= 4048;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 104;
        test_state <= test_b1_S4065;
      end
      test_b1_S4065: begin
        IMAGE_addr <= 4049;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 64;
        test_state <= test_b1_S4066;
      end
      test_b1_S4066: begin
        IMAGE_addr <= 4050;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 62;
        test_state <= test_b1_S4067;
      end
      test_b1_S4067: begin
        IMAGE_addr <= 4051;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4068;
      end
      test_b1_S4068: begin
        IMAGE_addr <= 4052;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4069;
      end
      test_b1_S4069: begin
        IMAGE_addr <= 4053;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4070;
      end
      test_b1_S4070: begin
        IMAGE_addr <= 4054;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S4071;
      end
      test_b1_S4071: begin
        IMAGE_addr <= 4055;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4072;
      end
      test_b1_S4072: begin
        IMAGE_addr <= 4056;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4073;
      end
      test_b1_S4073: begin
        IMAGE_addr <= 4057;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4041;
        test_state <= test_b1_S4074;
      end
      test_b1_S4074: begin
        IMAGE_addr <= 4058;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S4075;
      end
      test_b1_S4075: begin
        IMAGE_addr <= 4059;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4066;
        test_state <= test_b1_S4076;
      end
      test_b1_S4076: begin
        IMAGE_addr <= 4060;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S4077;
      end
      test_b1_S4077: begin
        IMAGE_addr <= 4061;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S4078;
      end
      test_b1_S4078: begin
        IMAGE_addr <= 4062;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 99;
        test_state <= test_b1_S4079;
      end
      test_b1_S4079: begin
        IMAGE_addr <= 4063;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 104;
        test_state <= test_b1_S4080;
      end
      test_b1_S4080: begin
        IMAGE_addr <= 4064;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 64;
        test_state <= test_b1_S4081;
      end
      test_b1_S4081: begin
        IMAGE_addr <= 4065;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4082;
      end
      test_b1_S4082: begin
        IMAGE_addr <= 4066;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4083;
      end
      test_b1_S4083: begin
        IMAGE_addr <= 4067;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4084;
      end
      test_b1_S4084: begin
        IMAGE_addr <= 4068;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S4085;
      end
      test_b1_S4085: begin
        IMAGE_addr <= 4069;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4074;
        test_state <= test_b1_S4086;
      end
      test_b1_S4086: begin
        IMAGE_addr <= 4070;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S4087;
      end
      test_b1_S4087: begin
        IMAGE_addr <= 4071;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4088;
      end
      test_b1_S4088: begin
        IMAGE_addr <= 4072;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 790;
        test_state <= test_b1_S4089;
      end
      test_b1_S4089: begin
        IMAGE_addr <= 4073;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4090;
      end
      test_b1_S4090: begin
        IMAGE_addr <= 4074;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S4091;
      end
      test_b1_S4091: begin
        IMAGE_addr <= 4075;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4078;
        test_state <= test_b1_S4092;
      end
      test_b1_S4092: begin
        IMAGE_addr <= 4076;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3978;
        test_state <= test_b1_S4093;
      end
      test_b1_S4093: begin
        IMAGE_addr <= 4077;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4094;
      end
      test_b1_S4094: begin
        IMAGE_addr <= 4078;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3735;
        test_state <= test_b1_S4095;
      end
      test_b1_S4095: begin
        IMAGE_addr <= 4079;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S4096;
      end
      test_b1_S4096: begin
        IMAGE_addr <= 4080;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4085;
        test_state <= test_b1_S4097;
      end
      test_b1_S4097: begin
        IMAGE_addr <= 4081;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S4098;
      end
      test_b1_S4098: begin
        IMAGE_addr <= 4082;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S4099;
      end
      test_b1_S4099: begin
        IMAGE_addr <= 4083;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 790;
        test_state <= test_b1_S4100;
      end
      test_b1_S4100: begin
        IMAGE_addr <= 4084;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4101;
      end
      test_b1_S4101: begin
        IMAGE_addr <= 4085;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S4102;
      end
      test_b1_S4102: begin
        IMAGE_addr <= 4086;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4089;
        test_state <= test_b1_S4103;
      end
      test_b1_S4103: begin
        IMAGE_addr <= 4087;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4006;
        test_state <= test_b1_S4104;
      end
      test_b1_S4104: begin
        IMAGE_addr <= 4088;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4105;
      end
      test_b1_S4105: begin
        IMAGE_addr <= 4089;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3735;
        test_state <= test_b1_S4106;
      end
      test_b1_S4106: begin
        IMAGE_addr <= 4090;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S4107;
      end
      test_b1_S4107: begin
        IMAGE_addr <= 4091;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4096;
        test_state <= test_b1_S4108;
      end
      test_b1_S4108: begin
        IMAGE_addr <= 4092;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S4109;
      end
      test_b1_S4109: begin
        IMAGE_addr <= 4093;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S4110;
      end
      test_b1_S4110: begin
        IMAGE_addr <= 4094;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 790;
        test_state <= test_b1_S4111;
      end
      test_b1_S4111: begin
        IMAGE_addr <= 4095;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4112;
      end
      test_b1_S4112: begin
        IMAGE_addr <= 4096;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S4113;
      end
      test_b1_S4113: begin
        IMAGE_addr <= 4097;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4103;
        test_state <= test_b1_S4114;
      end
      test_b1_S4114: begin
        IMAGE_addr <= 4098;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S4115;
      end
      test_b1_S4115: begin
        IMAGE_addr <= 4099;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 886;
        test_state <= test_b1_S4116;
      end
      test_b1_S4116: begin
        IMAGE_addr <= 4100;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 766;
        test_state <= test_b1_S4117;
      end
      test_b1_S4117: begin
        IMAGE_addr <= 4101;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4006;
        test_state <= test_b1_S4118;
      end
      test_b1_S4118: begin
        IMAGE_addr <= 4102;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4119;
      end
      test_b1_S4119: begin
        IMAGE_addr <= 4103;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3735;
        test_state <= test_b1_S4120;
      end
      test_b1_S4120: begin
        IMAGE_addr <= 4104;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S4121;
      end
      test_b1_S4121: begin
        IMAGE_addr <= 4105;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4110;
        test_state <= test_b1_S4122;
      end
      test_b1_S4122: begin
        IMAGE_addr <= 4106;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S4123;
      end
      test_b1_S4123: begin
        IMAGE_addr <= 4107;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S4124;
      end
      test_b1_S4124: begin
        IMAGE_addr <= 4108;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 790;
        test_state <= test_b1_S4125;
      end
      test_b1_S4125: begin
        IMAGE_addr <= 4109;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4126;
      end
      test_b1_S4126: begin
        IMAGE_addr <= 4110;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S4127;
      end
      test_b1_S4127: begin
        IMAGE_addr <= 4111;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4114;
        test_state <= test_b1_S4128;
      end
      test_b1_S4128: begin
        IMAGE_addr <= 4112;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4019;
        test_state <= test_b1_S4129;
      end
      test_b1_S4129: begin
        IMAGE_addr <= 4113;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4130;
      end
      test_b1_S4130: begin
        IMAGE_addr <= 4114;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3735;
        test_state <= test_b1_S4131;
      end
      test_b1_S4131: begin
        IMAGE_addr <= 4115;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4052;
        test_state <= test_b1_S4132;
      end
      test_b1_S4132: begin
        IMAGE_addr <= 4116;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4133;
      end
      test_b1_S4133: begin
        IMAGE_addr <= 4117;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4134;
      end
      test_b1_S4134: begin
        IMAGE_addr <= 4118;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4057;
        test_state <= test_b1_S4135;
      end
      test_b1_S4135: begin
        IMAGE_addr <= 4119;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S4136;
      end
      test_b1_S4136: begin
        IMAGE_addr <= 4120;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4126;
        test_state <= test_b1_S4137;
      end
      test_b1_S4137: begin
        IMAGE_addr <= 4121;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 99;
        test_state <= test_b1_S4138;
      end
      test_b1_S4138: begin
        IMAGE_addr <= 4122;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 111;
        test_state <= test_b1_S4139;
      end
      test_b1_S4139: begin
        IMAGE_addr <= 4123;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 112;
        test_state <= test_b1_S4140;
      end
      test_b1_S4140: begin
        IMAGE_addr <= 4124;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 121;
        test_state <= test_b1_S4141;
      end
      test_b1_S4141: begin
        IMAGE_addr <= 4125;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4142;
      end
      test_b1_S4142: begin
        IMAGE_addr <= 4126;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4143;
      end
      test_b1_S4143: begin
        IMAGE_addr <= 4127;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4144;
      end
      test_b1_S4144: begin
        IMAGE_addr <= 4128;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S4145;
      end
      test_b1_S4145: begin
        IMAGE_addr <= 4129;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4135;
        test_state <= test_b1_S4146;
      end
      test_b1_S4146: begin
        IMAGE_addr <= 4130;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S4147;
      end
      test_b1_S4147: begin
        IMAGE_addr <= 4131;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 189;
        test_state <= test_b1_S4148;
      end
      test_b1_S4148: begin
        IMAGE_addr <= 4132;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 766;
        test_state <= test_b1_S4149;
      end
      test_b1_S4149: begin
        IMAGE_addr <= 4133;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 197;
        test_state <= test_b1_S4150;
      end
      test_b1_S4150: begin
        IMAGE_addr <= 4134;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4151;
      end
      test_b1_S4151: begin
        IMAGE_addr <= 4135;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3841;
        test_state <= test_b1_S4152;
      end
      test_b1_S4152: begin
        IMAGE_addr <= 4136;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S4153;
      end
      test_b1_S4153: begin
        IMAGE_addr <= 4137;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S4154;
      end
      test_b1_S4154: begin
        IMAGE_addr <= 4138;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4155;
      end
      test_b1_S4155: begin
        IMAGE_addr <= 4139;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4156;
      end
      test_b1_S4156: begin
        IMAGE_addr <= 4140;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4118;
        test_state <= test_b1_S4157;
      end
      test_b1_S4157: begin
        IMAGE_addr <= 4141;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S4158;
      end
      test_b1_S4158: begin
        IMAGE_addr <= 4142;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4148;
        test_state <= test_b1_S4159;
      end
      test_b1_S4159: begin
        IMAGE_addr <= 4143;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 102;
        test_state <= test_b1_S4160;
      end
      test_b1_S4160: begin
        IMAGE_addr <= 4144;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S4161;
      end
      test_b1_S4161: begin
        IMAGE_addr <= 4145;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 108;
        test_state <= test_b1_S4162;
      end
      test_b1_S4162: begin
        IMAGE_addr <= 4146;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 108;
        test_state <= test_b1_S4163;
      end
      test_b1_S4163: begin
        IMAGE_addr <= 4147;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4164;
      end
      test_b1_S4164: begin
        IMAGE_addr <= 4148;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4165;
      end
      test_b1_S4165: begin
        IMAGE_addr <= 4149;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4166;
      end
      test_b1_S4166: begin
        IMAGE_addr <= 4150;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S4167;
      end
      test_b1_S4167: begin
        IMAGE_addr <= 4151;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 206;
        test_state <= test_b1_S4168;
      end
      test_b1_S4168: begin
        IMAGE_addr <= 4152;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S4169;
      end
      test_b1_S4169: begin
        IMAGE_addr <= 4153;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S4170;
      end
      test_b1_S4170: begin
        IMAGE_addr <= 4154;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4160;
        test_state <= test_b1_S4171;
      end
      test_b1_S4171: begin
        IMAGE_addr <= 4155;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 206;
        test_state <= test_b1_S4172;
      end
      test_b1_S4172: begin
        IMAGE_addr <= 4156;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S4173;
      end
      test_b1_S4173: begin
        IMAGE_addr <= 4157;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S4174;
      end
      test_b1_S4174: begin
        IMAGE_addr <= 4158;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 197;
        test_state <= test_b1_S4175;
      end
      test_b1_S4175: begin
        IMAGE_addr <= 4159;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4176;
      end
      test_b1_S4176: begin
        IMAGE_addr <= 4160;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3841;
        test_state <= test_b1_S4177;
      end
      test_b1_S4177: begin
        IMAGE_addr <= 4161;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S4178;
      end
      test_b1_S4178: begin
        IMAGE_addr <= 4162;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4179;
      end
      test_b1_S4179: begin
        IMAGE_addr <= 4163;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4180;
      end
      test_b1_S4180: begin
        IMAGE_addr <= 4164;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4140;
        test_state <= test_b1_S4181;
      end
      test_b1_S4181: begin
        IMAGE_addr <= 4165;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S4182;
      end
      test_b1_S4182: begin
        IMAGE_addr <= 4166;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4173;
        test_state <= test_b1_S4183;
      end
      test_b1_S4183: begin
        IMAGE_addr <= 4167;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S4184;
      end
      test_b1_S4184: begin
        IMAGE_addr <= 4168;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 104;
        test_state <= test_b1_S4185;
      end
      test_b1_S4185: begin
        IMAGE_addr <= 4169;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S4186;
      end
      test_b1_S4186: begin
        IMAGE_addr <= 4170;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S4187;
      end
      test_b1_S4187: begin
        IMAGE_addr <= 4171;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 100;
        test_state <= test_b1_S4188;
      end
      test_b1_S4188: begin
        IMAGE_addr <= 4172;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4189;
      end
      test_b1_S4189: begin
        IMAGE_addr <= 4173;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4190;
      end
      test_b1_S4190: begin
        IMAGE_addr <= 4174;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4191;
      end
      test_b1_S4191: begin
        IMAGE_addr <= 4175;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S4192;
      end
      test_b1_S4192: begin
        IMAGE_addr <= 4176;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8;
        test_state <= test_b1_S4193;
      end
      test_b1_S4193: begin
        IMAGE_addr <= 4177;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 213;
        test_state <= test_b1_S4194;
      end
      test_b1_S4194: begin
        IMAGE_addr <= 4178;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 206;
        test_state <= test_b1_S4195;
      end
      test_b1_S4195: begin
        IMAGE_addr <= 4179;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S4196;
      end
      test_b1_S4196: begin
        IMAGE_addr <= 4180;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4197;
      end
      test_b1_S4197: begin
        IMAGE_addr <= 4181;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 213;
        test_state <= test_b1_S4198;
      end
      test_b1_S4198: begin
        IMAGE_addr <= 4182;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4199;
      end
      test_b1_S4199: begin
        IMAGE_addr <= 4183;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4200;
      end
      test_b1_S4200: begin
        IMAGE_addr <= 4184;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4164;
        test_state <= test_b1_S4201;
      end
      test_b1_S4201: begin
        IMAGE_addr <= 4185;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3283;
        test_state <= test_b1_S4202;
      end
      test_b1_S4202: begin
        IMAGE_addr <= 4186;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4191;
        test_state <= test_b1_S4203;
      end
      test_b1_S4203: begin
        IMAGE_addr <= 4187;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S4204;
      end
      test_b1_S4204: begin
        IMAGE_addr <= 4188;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 102;
        test_state <= test_b1_S4205;
      end
      test_b1_S4205: begin
        IMAGE_addr <= 4189;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 59;
        test_state <= test_b1_S4206;
      end
      test_b1_S4206: begin
        IMAGE_addr <= 4190;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4207;
      end
      test_b1_S4207: begin
        IMAGE_addr <= 4191;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4208;
      end
      test_b1_S4208: begin
        IMAGE_addr <= 4192;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4209;
      end
      test_b1_S4209: begin
        IMAGE_addr <= 4193;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S4210;
      end
      test_b1_S4210: begin
        IMAGE_addr <= 4194;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 140;
        test_state <= test_b1_S4211;
      end
      test_b1_S4211: begin
        IMAGE_addr <= 4195;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S4212;
      end
      test_b1_S4212: begin
        IMAGE_addr <= 4196;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S4213;
      end
      test_b1_S4213: begin
        IMAGE_addr <= 4197;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 266;
        test_state <= test_b1_S4214;
      end
      test_b1_S4214: begin
        IMAGE_addr <= 4198;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3283;
        test_state <= test_b1_S4215;
      end
      test_b1_S4215: begin
        IMAGE_addr <= 4199;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S4216;
      end
      test_b1_S4216: begin
        IMAGE_addr <= 4200;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 52;
        test_state <= test_b1_S4217;
      end
      test_b1_S4217: begin
        IMAGE_addr <= 4201;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 323;
        test_state <= test_b1_S4218;
      end
      test_b1_S4218: begin
        IMAGE_addr <= 4202;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4219;
      end
      test_b1_S4219: begin
        IMAGE_addr <= 4203;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4220;
      end
      test_b1_S4220: begin
        IMAGE_addr <= 4204;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4184;
        test_state <= test_b1_S4221;
      end
      test_b1_S4221: begin
        IMAGE_addr <= 4205;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S4222;
      end
      test_b1_S4222: begin
        IMAGE_addr <= 4206;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4214;
        test_state <= test_b1_S4223;
      end
      test_b1_S4223: begin
        IMAGE_addr <= 4207;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 119;
        test_state <= test_b1_S4224;
      end
      test_b1_S4224: begin
        IMAGE_addr <= 4208;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S4225;
      end
      test_b1_S4225: begin
        IMAGE_addr <= 4209;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S4226;
      end
      test_b1_S4226: begin
        IMAGE_addr <= 4210;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 104;
        test_state <= test_b1_S4227;
      end
      test_b1_S4227: begin
        IMAGE_addr <= 4211;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S4228;
      end
      test_b1_S4228: begin
        IMAGE_addr <= 4212;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 110;
        test_state <= test_b1_S4229;
      end
      test_b1_S4229: begin
        IMAGE_addr <= 4213;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4230;
      end
      test_b1_S4230: begin
        IMAGE_addr <= 4214;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4231;
      end
      test_b1_S4231: begin
        IMAGE_addr <= 4215;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4232;
      end
      test_b1_S4232: begin
        IMAGE_addr <= 4216;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S4233;
      end
      test_b1_S4233: begin
        IMAGE_addr <= 4217;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 132;
        test_state <= test_b1_S4234;
      end
      test_b1_S4234: begin
        IMAGE_addr <= 4218;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 766;
        test_state <= test_b1_S4235;
      end
      test_b1_S4235: begin
        IMAGE_addr <= 4219;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 814;
        test_state <= test_b1_S4236;
      end
      test_b1_S4236: begin
        IMAGE_addr <= 4220;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S4237;
      end
      test_b1_S4237: begin
        IMAGE_addr <= 4221;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 806;
        test_state <= test_b1_S4238;
      end
      test_b1_S4238: begin
        IMAGE_addr <= 4222;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 766;
        test_state <= test_b1_S4239;
      end
      test_b1_S4239: begin
        IMAGE_addr <= 4223;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 20;
        test_state <= test_b1_S4240;
      end
      test_b1_S4240: begin
        IMAGE_addr <= 4224;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4241;
      end
      test_b1_S4241: begin
        IMAGE_addr <= 4225;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4242;
      end
      test_b1_S4242: begin
        IMAGE_addr <= 4226;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4204;
        test_state <= test_b1_S4243;
      end
      test_b1_S4243: begin
        IMAGE_addr <= 4227;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S4244;
      end
      test_b1_S4244: begin
        IMAGE_addr <= 4228;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4239;
        test_state <= test_b1_S4245;
      end
      test_b1_S4245: begin
        IMAGE_addr <= 4229;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 118;
        test_state <= test_b1_S4246;
      end
      test_b1_S4246: begin
        IMAGE_addr <= 4230;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S4247;
      end
      test_b1_S4247: begin
        IMAGE_addr <= 4231;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S4248;
      end
      test_b1_S4248: begin
        IMAGE_addr <= 4232;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S4249;
      end
      test_b1_S4249: begin
        IMAGE_addr <= 4233;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S4250;
      end
      test_b1_S4250: begin
        IMAGE_addr <= 4234;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 98;
        test_state <= test_b1_S4251;
      end
      test_b1_S4251: begin
        IMAGE_addr <= 4235;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 108;
        test_state <= test_b1_S4252;
      end
      test_b1_S4252: begin
        IMAGE_addr <= 4236;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S4253;
      end
      test_b1_S4253: begin
        IMAGE_addr <= 4237;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 58;
        test_state <= test_b1_S4254;
      end
      test_b1_S4254: begin
        IMAGE_addr <= 4238;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4255;
      end
      test_b1_S4255: begin
        IMAGE_addr <= 4239;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4256;
      end
      test_b1_S4256: begin
        IMAGE_addr <= 4240;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4257;
      end
      test_b1_S4257: begin
        IMAGE_addr <= 4241;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 621;
        test_state <= test_b1_S4258;
      end
      test_b1_S4258: begin
        IMAGE_addr <= 4242;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 213;
        test_state <= test_b1_S4259;
      end
      test_b1_S4259: begin
        IMAGE_addr <= 4243;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4260;
      end
      test_b1_S4260: begin
        IMAGE_addr <= 4244;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4261;
      end
      test_b1_S4261: begin
        IMAGE_addr <= 4245;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4226;
        test_state <= test_b1_S4262;
      end
      test_b1_S4262: begin
        IMAGE_addr <= 4246;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S4263;
      end
      test_b1_S4263: begin
        IMAGE_addr <= 4247;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4257;
        test_state <= test_b1_S4264;
      end
      test_b1_S4264: begin
        IMAGE_addr <= 4248;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 118;
        test_state <= test_b1_S4265;
      end
      test_b1_S4265: begin
        IMAGE_addr <= 4249;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S4266;
      end
      test_b1_S4266: begin
        IMAGE_addr <= 4250;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S4267;
      end
      test_b1_S4267: begin
        IMAGE_addr <= 4251;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S4268;
      end
      test_b1_S4268: begin
        IMAGE_addr <= 4252;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S4269;
      end
      test_b1_S4269: begin
        IMAGE_addr <= 4253;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 98;
        test_state <= test_b1_S4270;
      end
      test_b1_S4270: begin
        IMAGE_addr <= 4254;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 108;
        test_state <= test_b1_S4271;
      end
      test_b1_S4271: begin
        IMAGE_addr <= 4255;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S4272;
      end
      test_b1_S4272: begin
        IMAGE_addr <= 4256;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4273;
      end
      test_b1_S4273: begin
        IMAGE_addr <= 4257;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4274;
      end
      test_b1_S4274: begin
        IMAGE_addr <= 4258;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4275;
      end
      test_b1_S4275: begin
        IMAGE_addr <= 4259;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S4276;
      end
      test_b1_S4276: begin
        IMAGE_addr <= 4260;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4277;
      end
      test_b1_S4277: begin
        IMAGE_addr <= 4261;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4239;
        test_state <= test_b1_S4278;
      end
      test_b1_S4278: begin
        IMAGE_addr <= 4262;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4279;
      end
      test_b1_S4279: begin
        IMAGE_addr <= 4263;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4280;
      end
      test_b1_S4280: begin
        IMAGE_addr <= 4264;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4245;
        test_state <= test_b1_S4281;
      end
      test_b1_S4281: begin
        IMAGE_addr <= 4265;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S4282;
      end
      test_b1_S4282: begin
        IMAGE_addr <= 4266;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4276;
        test_state <= test_b1_S4283;
      end
      test_b1_S4283: begin
        IMAGE_addr <= 4267;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 99;
        test_state <= test_b1_S4284;
      end
      test_b1_S4284: begin
        IMAGE_addr <= 4268;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 111;
        test_state <= test_b1_S4285;
      end
      test_b1_S4285: begin
        IMAGE_addr <= 4269;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 110;
        test_state <= test_b1_S4286;
      end
      test_b1_S4286: begin
        IMAGE_addr <= 4270;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S4287;
      end
      test_b1_S4287: begin
        IMAGE_addr <= 4271;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S4288;
      end
      test_b1_S4288: begin
        IMAGE_addr <= 4272;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S4289;
      end
      test_b1_S4289: begin
        IMAGE_addr <= 4273;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 110;
        test_state <= test_b1_S4290;
      end
      test_b1_S4290: begin
        IMAGE_addr <= 4274;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S4291;
      end
      test_b1_S4291: begin
        IMAGE_addr <= 4275;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4292;
      end
      test_b1_S4292: begin
        IMAGE_addr <= 4276;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4293;
      end
      test_b1_S4293: begin
        IMAGE_addr <= 4277;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4294;
      end
      test_b1_S4294: begin
        IMAGE_addr <= 4278;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 621;
        test_state <= test_b1_S4295;
      end
      test_b1_S4295: begin
        IMAGE_addr <= 4279;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S4296;
      end
      test_b1_S4296: begin
        IMAGE_addr <= 4280;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S4297;
      end
      test_b1_S4297: begin
        IMAGE_addr <= 4281;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S4298;
      end
      test_b1_S4298: begin
        IMAGE_addr <= 4282;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 583;
        test_state <= test_b1_S4299;
      end
      test_b1_S4299: begin
        IMAGE_addr <= 4283;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S4300;
      end
      test_b1_S4300: begin
        IMAGE_addr <= 4284;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4301;
      end
      test_b1_S4301: begin
        IMAGE_addr <= 4285;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4302;
      end
      test_b1_S4302: begin
        IMAGE_addr <= 4286;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4264;
        test_state <= test_b1_S4303;
      end
      test_b1_S4303: begin
        IMAGE_addr <= 4287;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S4304;
      end
      test_b1_S4304: begin
        IMAGE_addr <= 4288;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4296;
        test_state <= test_b1_S4305;
      end
      test_b1_S4305: begin
        IMAGE_addr <= 4289;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S4306;
      end
      test_b1_S4306: begin
        IMAGE_addr <= 4290;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S4307;
      end
      test_b1_S4307: begin
        IMAGE_addr <= 4291;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S4308;
      end
      test_b1_S4308: begin
        IMAGE_addr <= 4292;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S4309;
      end
      test_b1_S4309: begin
        IMAGE_addr <= 4293;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 110;
        test_state <= test_b1_S4310;
      end
      test_b1_S4310: begin
        IMAGE_addr <= 4294;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 103;
        test_state <= test_b1_S4311;
      end
      test_b1_S4311: begin
        IMAGE_addr <= 4295;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4312;
      end
      test_b1_S4312: begin
        IMAGE_addr <= 4296;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4313;
      end
      test_b1_S4313: begin
        IMAGE_addr <= 4297;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4314;
      end
      test_b1_S4314: begin
        IMAGE_addr <= 4298;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 892;
        test_state <= test_b1_S4315;
      end
      test_b1_S4315: begin
        IMAGE_addr <= 4299;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4276;
        test_state <= test_b1_S4316;
      end
      test_b1_S4316: begin
        IMAGE_addr <= 4300;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4317;
      end
      test_b1_S4317: begin
        IMAGE_addr <= 4301;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4318;
      end
      test_b1_S4318: begin
        IMAGE_addr <= 4302;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4286;
        test_state <= test_b1_S4319;
      end
      test_b1_S4319: begin
        IMAGE_addr <= 4303;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S4320;
      end
      test_b1_S4320: begin
        IMAGE_addr <= 4304;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4311;
        test_state <= test_b1_S4321;
      end
      test_b1_S4321: begin
        IMAGE_addr <= 4305;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S4322;
      end
      test_b1_S4322: begin
        IMAGE_addr <= 4306;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 108;
        test_state <= test_b1_S4323;
      end
      test_b1_S4323: begin
        IMAGE_addr <= 4307;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 108;
        test_state <= test_b1_S4324;
      end
      test_b1_S4324: begin
        IMAGE_addr <= 4308;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 111;
        test_state <= test_b1_S4325;
      end
      test_b1_S4325: begin
        IMAGE_addr <= 4309;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S4326;
      end
      test_b1_S4326: begin
        IMAGE_addr <= 4310;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4327;
      end
      test_b1_S4327: begin
        IMAGE_addr <= 4311;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4328;
      end
      test_b1_S4328: begin
        IMAGE_addr <= 4312;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4329;
      end
      test_b1_S4329: begin
        IMAGE_addr <= 4313;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S4330;
      end
      test_b1_S4330: begin
        IMAGE_addr <= 4314;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S4331;
      end
      test_b1_S4331: begin
        IMAGE_addr <= 4315;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4332;
      end
      test_b1_S4332: begin
        IMAGE_addr <= 4316;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 822;
        test_state <= test_b1_S4333;
      end
      test_b1_S4333: begin
        IMAGE_addr <= 4317;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S4334;
      end
      test_b1_S4334: begin
        IMAGE_addr <= 4318;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4323;
        test_state <= test_b1_S4335;
      end
      test_b1_S4335: begin
        IMAGE_addr <= 4319;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S4336;
      end
      test_b1_S4336: begin
        IMAGE_addr <= 4320;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S4337;
      end
      test_b1_S4337: begin
        IMAGE_addr <= 4321;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2618;
        test_state <= test_b1_S4338;
      end
      test_b1_S4338: begin
        IMAGE_addr <= 4322;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4339;
      end
      test_b1_S4339: begin
        IMAGE_addr <= 4323;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S4340;
      end
      test_b1_S4340: begin
        IMAGE_addr <= 4324;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4333;
        test_state <= test_b1_S4341;
      end
      test_b1_S4341: begin
        IMAGE_addr <= 4325;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 25;
        test_state <= test_b1_S4342;
      end
      test_b1_S4342: begin
        IMAGE_addr <= 4326;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 27;
        test_state <= test_b1_S4343;
      end
      test_b1_S4343: begin
        IMAGE_addr <= 4327;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S4344;
      end
      test_b1_S4344: begin
        IMAGE_addr <= 4328;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4345;
      end
      test_b1_S4345: begin
        IMAGE_addr <= 4329;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 213;
        test_state <= test_b1_S4346;
      end
      test_b1_S4346: begin
        IMAGE_addr <= 4330;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8;
        test_state <= test_b1_S4347;
      end
      test_b1_S4347: begin
        IMAGE_addr <= 4331;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4325;
        test_state <= test_b1_S4348;
      end
      test_b1_S4348: begin
        IMAGE_addr <= 4332;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4349;
      end
      test_b1_S4349: begin
        IMAGE_addr <= 4333;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 732;
        test_state <= test_b1_S4350;
      end
      test_b1_S4350: begin
        IMAGE_addr <= 4334;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4351;
      end
      test_b1_S4351: begin
        IMAGE_addr <= 4335;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4352;
      end
      test_b1_S4352: begin
        IMAGE_addr <= 4336;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4302;
        test_state <= test_b1_S4353;
      end
      test_b1_S4353: begin
        IMAGE_addr <= 4337;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S4354;
      end
      test_b1_S4354: begin
        IMAGE_addr <= 4338;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4344;
        test_state <= test_b1_S4355;
      end
      test_b1_S4355: begin
        IMAGE_addr <= 4339;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 108;
        test_state <= test_b1_S4356;
      end
      test_b1_S4356: begin
        IMAGE_addr <= 4340;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S4357;
      end
      test_b1_S4357: begin
        IMAGE_addr <= 4341;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S4358;
      end
      test_b1_S4358: begin
        IMAGE_addr <= 4342;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S4359;
      end
      test_b1_S4359: begin
        IMAGE_addr <= 4343;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4360;
      end
      test_b1_S4360: begin
        IMAGE_addr <= 4344;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 206;
        test_state <= test_b1_S4361;
      end
      test_b1_S4361: begin
        IMAGE_addr <= 4345;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S4362;
      end
      test_b1_S4362: begin
        IMAGE_addr <= 4346;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4311;
        test_state <= test_b1_S4363;
      end
      test_b1_S4363: begin
        IMAGE_addr <= 4347;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4364;
      end
      test_b1_S4364: begin
        IMAGE_addr <= 4348;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4365;
      end
      test_b1_S4365: begin
        IMAGE_addr <= 4349;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4336;
        test_state <= test_b1_S4366;
      end
      test_b1_S4366: begin
        IMAGE_addr <= 4350;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S4367;
      end
      test_b1_S4367: begin
        IMAGE_addr <= 4351;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4360;
        test_state <= test_b1_S4368;
      end
      test_b1_S4368: begin
        IMAGE_addr <= 4352;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S4369;
      end
      test_b1_S4369: begin
        IMAGE_addr <= 4353;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 108;
        test_state <= test_b1_S4370;
      end
      test_b1_S4370: begin
        IMAGE_addr <= 4354;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S4371;
      end
      test_b1_S4371: begin
        IMAGE_addr <= 4355;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 109;
        test_state <= test_b1_S4372;
      end
      test_b1_S4372: begin
        IMAGE_addr <= 4356;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S4373;
      end
      test_b1_S4373: begin
        IMAGE_addr <= 4357;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 110;
        test_state <= test_b1_S4374;
      end
      test_b1_S4374: begin
        IMAGE_addr <= 4358;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S4375;
      end
      test_b1_S4375: begin
        IMAGE_addr <= 4359;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4376;
      end
      test_b1_S4376: begin
        IMAGE_addr <= 4360;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 621;
        test_state <= test_b1_S4377;
      end
      test_b1_S4377: begin
        IMAGE_addr <= 4361;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S4378;
      end
      test_b1_S4378: begin
        IMAGE_addr <= 4362;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S4379;
      end
      test_b1_S4379: begin
        IMAGE_addr <= 4363;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S4380;
      end
      test_b1_S4380: begin
        IMAGE_addr <= 4364;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S4381;
      end
      test_b1_S4381: begin
        IMAGE_addr <= 4365;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 583;
        test_state <= test_b1_S4382;
      end
      test_b1_S4382: begin
        IMAGE_addr <= 4366;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S4383;
      end
      test_b1_S4383: begin
        IMAGE_addr <= 4367;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 26;
        test_state <= test_b1_S4384;
      end
      test_b1_S4384: begin
        IMAGE_addr <= 4368;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4385;
      end
      test_b1_S4385: begin
        IMAGE_addr <= 4369;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4386;
      end
      test_b1_S4386: begin
        IMAGE_addr <= 4370;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4302;
        test_state <= test_b1_S4387;
      end
      test_b1_S4387: begin
        IMAGE_addr <= 4371;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S4388;
      end
      test_b1_S4388: begin
        IMAGE_addr <= 4372;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4382;
        test_state <= test_b1_S4389;
      end
      test_b1_S4389: begin
        IMAGE_addr <= 4373;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S4390;
      end
      test_b1_S4390: begin
        IMAGE_addr <= 4374;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 108;
        test_state <= test_b1_S4391;
      end
      test_b1_S4391: begin
        IMAGE_addr <= 4375;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S4392;
      end
      test_b1_S4392: begin
        IMAGE_addr <= 4376;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 109;
        test_state <= test_b1_S4393;
      end
      test_b1_S4393: begin
        IMAGE_addr <= 4377;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S4394;
      end
      test_b1_S4394: begin
        IMAGE_addr <= 4378;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 110;
        test_state <= test_b1_S4395;
      end
      test_b1_S4395: begin
        IMAGE_addr <= 4379;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S4396;
      end
      test_b1_S4396: begin
        IMAGE_addr <= 4380;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S4397;
      end
      test_b1_S4397: begin
        IMAGE_addr <= 4381;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4398;
      end
      test_b1_S4398: begin
        IMAGE_addr <= 4382;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4399;
      end
      test_b1_S4399: begin
        IMAGE_addr <= 4383;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4400;
      end
      test_b1_S4400: begin
        IMAGE_addr <= 4384;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S4401;
      end
      test_b1_S4401: begin
        IMAGE_addr <= 4385;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4344;
        test_state <= test_b1_S4402;
      end
      test_b1_S4402: begin
        IMAGE_addr <= 4386;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S4403;
      end
      test_b1_S4403: begin
        IMAGE_addr <= 4387;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S4404;
      end
      test_b1_S4404: begin
        IMAGE_addr <= 4388;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4360;
        test_state <= test_b1_S4405;
      end
      test_b1_S4405: begin
        IMAGE_addr <= 4389;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3841;
        test_state <= test_b1_S4406;
      end
      test_b1_S4406: begin
        IMAGE_addr <= 4390;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S4407;
      end
      test_b1_S4407: begin
        IMAGE_addr <= 4391;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4408;
      end
      test_b1_S4408: begin
        IMAGE_addr <= 4392;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4409;
      end
      test_b1_S4409: begin
        IMAGE_addr <= 4393;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4370;
        test_state <= test_b1_S4410;
      end
      test_b1_S4410: begin
        IMAGE_addr <= 4394;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S4411;
      end
      test_b1_S4411: begin
        IMAGE_addr <= 4395;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4404;
        test_state <= test_b1_S4412;
      end
      test_b1_S4412: begin
        IMAGE_addr <= 4396;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 100;
        test_state <= test_b1_S4413;
      end
      test_b1_S4413: begin
        IMAGE_addr <= 4397;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S4414;
      end
      test_b1_S4414: begin
        IMAGE_addr <= 4398;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 99;
        test_state <= test_b1_S4415;
      end
      test_b1_S4415: begin
        IMAGE_addr <= 4399;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S4416;
      end
      test_b1_S4416: begin
        IMAGE_addr <= 4400;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 109;
        test_state <= test_b1_S4417;
      end
      test_b1_S4417: begin
        IMAGE_addr <= 4401;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S4418;
      end
      test_b1_S4418: begin
        IMAGE_addr <= 4402;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 108;
        test_state <= test_b1_S4419;
      end
      test_b1_S4419: begin
        IMAGE_addr <= 4403;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4420;
      end
      test_b1_S4420: begin
        IMAGE_addr <= 4404;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4421;
      end
      test_b1_S4421: begin
        IMAGE_addr <= 4405;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4422;
      end
      test_b1_S4422: begin
        IMAGE_addr <= 4406;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S4423;
      end
      test_b1_S4423: begin
        IMAGE_addr <= 4407;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 10;
        test_state <= test_b1_S4424;
      end
      test_b1_S4424: begin
        IMAGE_addr <= 4408;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S4425;
      end
      test_b1_S4425: begin
        IMAGE_addr <= 4409;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 925;
        test_state <= test_b1_S4426;
      end
      test_b1_S4426: begin
        IMAGE_addr <= 4410;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S4427;
      end
      test_b1_S4427: begin
        IMAGE_addr <= 4411;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4428;
      end
      test_b1_S4428: begin
        IMAGE_addr <= 4412;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4429;
      end
      test_b1_S4429: begin
        IMAGE_addr <= 4413;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4393;
        test_state <= test_b1_S4430;
      end
      test_b1_S4430: begin
        IMAGE_addr <= 4414;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S4431;
      end
      test_b1_S4431: begin
        IMAGE_addr <= 4415;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4420;
        test_state <= test_b1_S4432;
      end
      test_b1_S4432: begin
        IMAGE_addr <= 4416;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 104;
        test_state <= test_b1_S4433;
      end
      test_b1_S4433: begin
        IMAGE_addr <= 4417;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S4434;
      end
      test_b1_S4434: begin
        IMAGE_addr <= 4418;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 120;
        test_state <= test_b1_S4435;
      end
      test_b1_S4435: begin
        IMAGE_addr <= 4419;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4436;
      end
      test_b1_S4436: begin
        IMAGE_addr <= 4420;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4437;
      end
      test_b1_S4437: begin
        IMAGE_addr <= 4421;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4438;
      end
      test_b1_S4438: begin
        IMAGE_addr <= 4422;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S4439;
      end
      test_b1_S4439: begin
        IMAGE_addr <= 4423;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 16;
        test_state <= test_b1_S4440;
      end
      test_b1_S4440: begin
        IMAGE_addr <= 4424;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S4441;
      end
      test_b1_S4441: begin
        IMAGE_addr <= 4425;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 925;
        test_state <= test_b1_S4442;
      end
      test_b1_S4442: begin
        IMAGE_addr <= 4426;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S4443;
      end
      test_b1_S4443: begin
        IMAGE_addr <= 4427;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4444;
      end
      test_b1_S4444: begin
        IMAGE_addr <= 4428;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4445;
      end
      test_b1_S4445: begin
        IMAGE_addr <= 4429;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4413;
        test_state <= test_b1_S4446;
      end
      test_b1_S4446: begin
        IMAGE_addr <= 4430;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S4447;
      end
      test_b1_S4447: begin
        IMAGE_addr <= 4431;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4438;
        test_state <= test_b1_S4448;
      end
      test_b1_S4448: begin
        IMAGE_addr <= 4432;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 111;
        test_state <= test_b1_S4449;
      end
      test_b1_S4449: begin
        IMAGE_addr <= 4433;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 99;
        test_state <= test_b1_S4450;
      end
      test_b1_S4450: begin
        IMAGE_addr <= 4434;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S4451;
      end
      test_b1_S4451: begin
        IMAGE_addr <= 4435;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S4452;
      end
      test_b1_S4452: begin
        IMAGE_addr <= 4436;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 108;
        test_state <= test_b1_S4453;
      end
      test_b1_S4453: begin
        IMAGE_addr <= 4437;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4454;
      end
      test_b1_S4454: begin
        IMAGE_addr <= 4438;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4455;
      end
      test_b1_S4455: begin
        IMAGE_addr <= 4439;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4456;
      end
      test_b1_S4456: begin
        IMAGE_addr <= 4440;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S4457;
      end
      test_b1_S4457: begin
        IMAGE_addr <= 4441;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8;
        test_state <= test_b1_S4458;
      end
      test_b1_S4458: begin
        IMAGE_addr <= 4442;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S4459;
      end
      test_b1_S4459: begin
        IMAGE_addr <= 4443;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 925;
        test_state <= test_b1_S4460;
      end
      test_b1_S4460: begin
        IMAGE_addr <= 4444;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S4461;
      end
      test_b1_S4461: begin
        IMAGE_addr <= 4445;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4462;
      end
      test_b1_S4462: begin
        IMAGE_addr <= 4446;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4463;
      end
      test_b1_S4463: begin
        IMAGE_addr <= 4447;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4429;
        test_state <= test_b1_S4464;
      end
      test_b1_S4464: begin
        IMAGE_addr <= 4448;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S4465;
      end
      test_b1_S4465: begin
        IMAGE_addr <= 4449;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4457;
        test_state <= test_b1_S4466;
      end
      test_b1_S4466: begin
        IMAGE_addr <= 4450;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 98;
        test_state <= test_b1_S4467;
      end
      test_b1_S4467: begin
        IMAGE_addr <= 4451;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S4468;
      end
      test_b1_S4468: begin
        IMAGE_addr <= 4452;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 110;
        test_state <= test_b1_S4469;
      end
      test_b1_S4469: begin
        IMAGE_addr <= 4453;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S4470;
      end
      test_b1_S4470: begin
        IMAGE_addr <= 4454;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S4471;
      end
      test_b1_S4471: begin
        IMAGE_addr <= 4455;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 121;
        test_state <= test_b1_S4472;
      end
      test_b1_S4472: begin
        IMAGE_addr <= 4456;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4473;
      end
      test_b1_S4473: begin
        IMAGE_addr <= 4457;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4474;
      end
      test_b1_S4474: begin
        IMAGE_addr <= 4458;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4475;
      end
      test_b1_S4475: begin
        IMAGE_addr <= 4459;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S4476;
      end
      test_b1_S4476: begin
        IMAGE_addr <= 4460;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S4477;
      end
      test_b1_S4477: begin
        IMAGE_addr <= 4461;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S4478;
      end
      test_b1_S4478: begin
        IMAGE_addr <= 4462;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 925;
        test_state <= test_b1_S4479;
      end
      test_b1_S4479: begin
        IMAGE_addr <= 4463;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S4480;
      end
      test_b1_S4480: begin
        IMAGE_addr <= 4464;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4481;
      end
      test_b1_S4481: begin
        IMAGE_addr <= 4465;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4482;
      end
      test_b1_S4482: begin
        IMAGE_addr <= 4466;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4447;
        test_state <= test_b1_S4483;
      end
      test_b1_S4483: begin
        IMAGE_addr <= 4467;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 310;
        test_state <= test_b1_S4484;
      end
      test_b1_S4484: begin
        IMAGE_addr <= 4468;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4473;
        test_state <= test_b1_S4485;
      end
      test_b1_S4485: begin
        IMAGE_addr <= 4469;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 98;
        test_state <= test_b1_S4486;
      end
      test_b1_S4486: begin
        IMAGE_addr <= 4470;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 117;
        test_state <= test_b1_S4487;
      end
      test_b1_S4487: begin
        IMAGE_addr <= 4471;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 102;
        test_state <= test_b1_S4488;
      end
      test_b1_S4488: begin
        IMAGE_addr <= 4472;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4489;
      end
      test_b1_S4489: begin
        IMAGE_addr <= 4473;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 48;
        test_state <= test_b1_S4490;
      end
      test_b1_S4490: begin
        IMAGE_addr <= 4474;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4491;
      end
      test_b1_S4491: begin
        IMAGE_addr <= 4475;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4492;
      end
      test_b1_S4492: begin
        IMAGE_addr <= 4476;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4493;
      end
      test_b1_S4493: begin
        IMAGE_addr <= 4477;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4494;
      end
      test_b1_S4494: begin
        IMAGE_addr <= 4478;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4495;
      end
      test_b1_S4495: begin
        IMAGE_addr <= 4479;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4496;
      end
      test_b1_S4496: begin
        IMAGE_addr <= 4480;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4497;
      end
      test_b1_S4497: begin
        IMAGE_addr <= 4481;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4498;
      end
      test_b1_S4498: begin
        IMAGE_addr <= 4482;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4499;
      end
      test_b1_S4499: begin
        IMAGE_addr <= 4483;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4500;
      end
      test_b1_S4500: begin
        IMAGE_addr <= 4484;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4501;
      end
      test_b1_S4501: begin
        IMAGE_addr <= 4485;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4502;
      end
      test_b1_S4502: begin
        IMAGE_addr <= 4486;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4503;
      end
      test_b1_S4503: begin
        IMAGE_addr <= 4487;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4504;
      end
      test_b1_S4504: begin
        IMAGE_addr <= 4488;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4505;
      end
      test_b1_S4505: begin
        IMAGE_addr <= 4489;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4506;
      end
      test_b1_S4506: begin
        IMAGE_addr <= 4490;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4507;
      end
      test_b1_S4507: begin
        IMAGE_addr <= 4491;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4508;
      end
      test_b1_S4508: begin
        IMAGE_addr <= 4492;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4509;
      end
      test_b1_S4509: begin
        IMAGE_addr <= 4493;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4510;
      end
      test_b1_S4510: begin
        IMAGE_addr <= 4494;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4511;
      end
      test_b1_S4511: begin
        IMAGE_addr <= 4495;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4512;
      end
      test_b1_S4512: begin
        IMAGE_addr <= 4496;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4513;
      end
      test_b1_S4513: begin
        IMAGE_addr <= 4497;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4514;
      end
      test_b1_S4514: begin
        IMAGE_addr <= 4498;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4515;
      end
      test_b1_S4515: begin
        IMAGE_addr <= 4499;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4516;
      end
      test_b1_S4516: begin
        IMAGE_addr <= 4500;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4517;
      end
      test_b1_S4517: begin
        IMAGE_addr <= 4501;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4518;
      end
      test_b1_S4518: begin
        IMAGE_addr <= 4502;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4519;
      end
      test_b1_S4519: begin
        IMAGE_addr <= 4503;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4520;
      end
      test_b1_S4520: begin
        IMAGE_addr <= 4504;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4521;
      end
      test_b1_S4521: begin
        IMAGE_addr <= 4505;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S4522;
      end
      test_b1_S4522: begin
        IMAGE_addr <= 4506;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4523;
      end
      test_b1_S4523: begin
        IMAGE_addr <= 4507;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4466;
        test_state <= test_b1_S4524;
      end
      test_b1_S4524: begin
        IMAGE_addr <= 4508;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 310;
        test_state <= test_b1_S4525;
      end
      test_b1_S4525: begin
        IMAGE_addr <= 4509;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4505;
        test_state <= test_b1_S4526;
      end
      test_b1_S4526: begin
        IMAGE_addr <= 4510;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 100;
        test_state <= test_b1_S4527;
      end
      test_b1_S4527: begin
        IMAGE_addr <= 4511;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S4528;
      end
      test_b1_S4528: begin
        IMAGE_addr <= 4512;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 103;
        test_state <= test_b1_S4529;
      end
      test_b1_S4529: begin
        IMAGE_addr <= 4513;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S4530;
      end
      test_b1_S4530: begin
        IMAGE_addr <= 4514;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S4531;
      end
      test_b1_S4531: begin
        IMAGE_addr <= 4515;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S4532;
      end
      test_b1_S4532: begin
        IMAGE_addr <= 4516;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4533;
      end
      test_b1_S4533: begin
        IMAGE_addr <= 4517;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4507;
        test_state <= test_b1_S4534;
      end
      test_b1_S4534: begin
        IMAGE_addr <= 4518;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 310;
        test_state <= test_b1_S4535;
      end
      test_b1_S4535: begin
        IMAGE_addr <= 4519;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4506;
        test_state <= test_b1_S4536;
      end
      test_b1_S4536: begin
        IMAGE_addr <= 4520;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 112;
        test_state <= test_b1_S4537;
      end
      test_b1_S4537: begin
        IMAGE_addr <= 4521;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 111;
        test_state <= test_b1_S4538;
      end
      test_b1_S4538: begin
        IMAGE_addr <= 4522;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S4539;
      end
      test_b1_S4539: begin
        IMAGE_addr <= 4523;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4540;
      end
      test_b1_S4540: begin
        IMAGE_addr <= 4524;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4517;
        test_state <= test_b1_S4541;
      end
      test_b1_S4541: begin
        IMAGE_addr <= 4525;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S4542;
      end
      test_b1_S4542: begin
        IMAGE_addr <= 4526;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4533;
        test_state <= test_b1_S4543;
      end
      test_b1_S4543: begin
        IMAGE_addr <= 4527;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S4544;
      end
      test_b1_S4544: begin
        IMAGE_addr <= 4528;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 112;
        test_state <= test_b1_S4545;
      end
      test_b1_S4545: begin
        IMAGE_addr <= 4529;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 108;
        test_state <= test_b1_S4546;
      end
      test_b1_S4546: begin
        IMAGE_addr <= 4530;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S4547;
      end
      test_b1_S4547: begin
        IMAGE_addr <= 4531;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S4548;
      end
      test_b1_S4548: begin
        IMAGE_addr <= 4532;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4549;
      end
      test_b1_S4549: begin
        IMAGE_addr <= 4533;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S4550;
      end
      test_b1_S4550: begin
        IMAGE_addr <= 4534;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 925;
        test_state <= test_b1_S4551;
      end
      test_b1_S4551: begin
        IMAGE_addr <= 4535;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S4552;
      end
      test_b1_S4552: begin
        IMAGE_addr <= 4536;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 19;
        test_state <= test_b1_S4553;
      end
      test_b1_S4553: begin
        IMAGE_addr <= 4537;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S4554;
      end
      test_b1_S4554: begin
        IMAGE_addr <= 4538;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 943;
        test_state <= test_b1_S4555;
      end
      test_b1_S4555: begin
        IMAGE_addr <= 4539;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 16;
        test_state <= test_b1_S4556;
      end
      test_b1_S4556: begin
        IMAGE_addr <= 4540;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S4557;
      end
      test_b1_S4557: begin
        IMAGE_addr <= 4541;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S4558;
      end
      test_b1_S4558: begin
        IMAGE_addr <= 4542;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S4559;
      end
      test_b1_S4559: begin
        IMAGE_addr <= 4543;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4505;
        test_state <= test_b1_S4560;
      end
      test_b1_S4560: begin
        IMAGE_addr <= 4544;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2651;
        test_state <= test_b1_S4561;
      end
      test_b1_S4561: begin
        IMAGE_addr <= 4545;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 25;
        test_state <= test_b1_S4562;
      end
      test_b1_S4562: begin
        IMAGE_addr <= 4546;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8;
        test_state <= test_b1_S4563;
      end
      test_b1_S4563: begin
        IMAGE_addr <= 4547;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4533;
        test_state <= test_b1_S4564;
      end
      test_b1_S4564: begin
        IMAGE_addr <= 4548;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4565;
      end
      test_b1_S4565: begin
        IMAGE_addr <= 4549;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4566;
      end
      test_b1_S4566: begin
        IMAGE_addr <= 4550;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4524;
        test_state <= test_b1_S4567;
      end
      test_b1_S4567: begin
        IMAGE_addr <= 4551;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S4568;
      end
      test_b1_S4568: begin
        IMAGE_addr <= 4552;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4559;
        test_state <= test_b1_S4569;
      end
      test_b1_S4569: begin
        IMAGE_addr <= 4553;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 98;
        test_state <= test_b1_S4570;
      end
      test_b1_S4570: begin
        IMAGE_addr <= 4554;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 117;
        test_state <= test_b1_S4571;
      end
      test_b1_S4571: begin
        IMAGE_addr <= 4555;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S4572;
      end
      test_b1_S4572: begin
        IMAGE_addr <= 4556;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 108;
        test_state <= test_b1_S4573;
      end
      test_b1_S4573: begin
        IMAGE_addr <= 4557;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 100;
        test_state <= test_b1_S4574;
      end
      test_b1_S4574: begin
        IMAGE_addr <= 4558;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4575;
      end
      test_b1_S4575: begin
        IMAGE_addr <= 4559;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S4576;
      end
      test_b1_S4576: begin
        IMAGE_addr <= 4560;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4473;
        test_state <= test_b1_S4577;
      end
      test_b1_S4577: begin
        IMAGE_addr <= 4561;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S4578;
      end
      test_b1_S4578: begin
        IMAGE_addr <= 4562;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4506;
        test_state <= test_b1_S4579;
      end
      test_b1_S4579: begin
        IMAGE_addr <= 4563;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S4580;
      end
      test_b1_S4580: begin
        IMAGE_addr <= 4564;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S4581;
      end
      test_b1_S4581: begin
        IMAGE_addr <= 4565;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4572;
        test_state <= test_b1_S4582;
      end
      test_b1_S4582: begin
        IMAGE_addr <= 4566;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S4583;
      end
      test_b1_S4583: begin
        IMAGE_addr <= 4567;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4506;
        test_state <= test_b1_S4584;
      end
      test_b1_S4584: begin
        IMAGE_addr <= 4568;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S4585;
      end
      test_b1_S4585: begin
        IMAGE_addr <= 4569;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S4586;
      end
      test_b1_S4586: begin
        IMAGE_addr <= 4570;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 197;
        test_state <= test_b1_S4587;
      end
      test_b1_S4587: begin
        IMAGE_addr <= 4571;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4588;
      end
      test_b1_S4588: begin
        IMAGE_addr <= 4572;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 751;
        test_state <= test_b1_S4589;
      end
      test_b1_S4589: begin
        IMAGE_addr <= 4573;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S4590;
      end
      test_b1_S4590: begin
        IMAGE_addr <= 4574;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4505;
        test_state <= test_b1_S4591;
      end
      test_b1_S4591: begin
        IMAGE_addr <= 4575;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S4592;
      end
      test_b1_S4592: begin
        IMAGE_addr <= 4576;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S4593;
      end
      test_b1_S4593: begin
        IMAGE_addr <= 4577;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4580;
        test_state <= test_b1_S4594;
      end
      test_b1_S4594: begin
        IMAGE_addr <= 4578;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 197;
        test_state <= test_b1_S4595;
      end
      test_b1_S4595: begin
        IMAGE_addr <= 4579;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4596;
      end
      test_b1_S4596: begin
        IMAGE_addr <= 4580;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3841;
        test_state <= test_b1_S4597;
      end
      test_b1_S4597: begin
        IMAGE_addr <= 4581;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S4598;
      end
      test_b1_S4598: begin
        IMAGE_addr <= 4582;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4599;
      end
      test_b1_S4599: begin
        IMAGE_addr <= 4583;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S4600;
      end
      test_b1_S4600: begin
        IMAGE_addr <= 4584;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S4601;
      end
      test_b1_S4601: begin
        IMAGE_addr <= 4585;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4602;
      end
      test_b1_S4602: begin
        IMAGE_addr <= 4586;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4603;
      end
      test_b1_S4603: begin
        IMAGE_addr <= 4587;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4550;
        test_state <= test_b1_S4604;
      end
      test_b1_S4604: begin
        IMAGE_addr <= 4588;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S4605;
      end
      test_b1_S4605: begin
        IMAGE_addr <= 4589;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4598;
        test_state <= test_b1_S4606;
      end
      test_b1_S4606: begin
        IMAGE_addr <= 4590;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 110;
        test_state <= test_b1_S4607;
      end
      test_b1_S4607: begin
        IMAGE_addr <= 4591;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S4608;
      end
      test_b1_S4608: begin
        IMAGE_addr <= 4592;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 103;
        test_state <= test_b1_S4609;
      end
      test_b1_S4609: begin
        IMAGE_addr <= 4593;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S4610;
      end
      test_b1_S4610: begin
        IMAGE_addr <= 4594;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S4611;
      end
      test_b1_S4611: begin
        IMAGE_addr <= 4595;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S4612;
      end
      test_b1_S4612: begin
        IMAGE_addr <= 4596;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 63;
        test_state <= test_b1_S4613;
      end
      test_b1_S4613: begin
        IMAGE_addr <= 4597;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4614;
      end
      test_b1_S4614: begin
        IMAGE_addr <= 4598;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S4615;
      end
      test_b1_S4615: begin
        IMAGE_addr <= 4599;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S4616;
      end
      test_b1_S4616: begin
        IMAGE_addr <= 4600;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4617;
      end
      test_b1_S4617: begin
        IMAGE_addr <= 4601;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 806;
        test_state <= test_b1_S4618;
      end
      test_b1_S4618: begin
        IMAGE_addr <= 4602;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 140;
        test_state <= test_b1_S4619;
      end
      test_b1_S4619: begin
        IMAGE_addr <= 4603;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 25;
        test_state <= test_b1_S4620;
      end
      test_b1_S4620: begin
        IMAGE_addr <= 4604;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S4621;
      end
      test_b1_S4621: begin
        IMAGE_addr <= 4605;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 176;
        test_state <= test_b1_S4622;
      end
      test_b1_S4622: begin
        IMAGE_addr <= 4606;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S4623;
      end
      test_b1_S4623: begin
        IMAGE_addr <= 4607;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 45;
        test_state <= test_b1_S4624;
      end
      test_b1_S4624: begin
        IMAGE_addr <= 4608;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S4625;
      end
      test_b1_S4625: begin
        IMAGE_addr <= 4609;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4506;
        test_state <= test_b1_S4626;
      end
      test_b1_S4626: begin
        IMAGE_addr <= 4610;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S4627;
      end
      test_b1_S4627: begin
        IMAGE_addr <= 4611;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4628;
      end
      test_b1_S4628: begin
        IMAGE_addr <= 4612;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4629;
      end
      test_b1_S4629: begin
        IMAGE_addr <= 4613;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4447;
        test_state <= test_b1_S4630;
      end
      test_b1_S4630: begin
        IMAGE_addr <= 4614;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S4631;
      end
      test_b1_S4631: begin
        IMAGE_addr <= 4615;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4625;
        test_state <= test_b1_S4632;
      end
      test_b1_S4632: begin
        IMAGE_addr <= 4616;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S4633;
      end
      test_b1_S4633: begin
        IMAGE_addr <= 4617;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 111;
        test_state <= test_b1_S4634;
      end
      test_b1_S4634: begin
        IMAGE_addr <= 4618;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 83;
        test_state <= test_b1_S4635;
      end
      test_b1_S4635: begin
        IMAGE_addr <= 4619;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S4636;
      end
      test_b1_S4636: begin
        IMAGE_addr <= 4620;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S4637;
      end
      test_b1_S4637: begin
        IMAGE_addr <= 4621;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S4638;
      end
      test_b1_S4638: begin
        IMAGE_addr <= 4622;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 110;
        test_state <= test_b1_S4639;
      end
      test_b1_S4639: begin
        IMAGE_addr <= 4623;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 103;
        test_state <= test_b1_S4640;
      end
      test_b1_S4640: begin
        IMAGE_addr <= 4624;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4641;
      end
      test_b1_S4641: begin
        IMAGE_addr <= 4625;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4642;
      end
      test_b1_S4642: begin
        IMAGE_addr <= 4626;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4643;
      end
      test_b1_S4643: begin
        IMAGE_addr <= 4627;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S4644;
      end
      test_b1_S4644: begin
        IMAGE_addr <= 4628;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4645;
      end
      test_b1_S4645: begin
        IMAGE_addr <= 4629;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S4646;
      end
      test_b1_S4646: begin
        IMAGE_addr <= 4630;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4635;
        test_state <= test_b1_S4647;
      end
      test_b1_S4647: begin
        IMAGE_addr <= 4631;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S4648;
      end
      test_b1_S4648: begin
        IMAGE_addr <= 4632;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4506;
        test_state <= test_b1_S4649;
      end
      test_b1_S4649: begin
        IMAGE_addr <= 4633;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S4650;
      end
      test_b1_S4650: begin
        IMAGE_addr <= 4634;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4651;
      end
      test_b1_S4651: begin
        IMAGE_addr <= 4635;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S4652;
      end
      test_b1_S4652: begin
        IMAGE_addr <= 4636;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4641;
        test_state <= test_b1_S4653;
      end
      test_b1_S4653: begin
        IMAGE_addr <= 4637;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S4654;
      end
      test_b1_S4654: begin
        IMAGE_addr <= 4638;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4505;
        test_state <= test_b1_S4655;
      end
      test_b1_S4655: begin
        IMAGE_addr <= 4639;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S4656;
      end
      test_b1_S4656: begin
        IMAGE_addr <= 4640;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4657;
      end
      test_b1_S4657: begin
        IMAGE_addr <= 4641;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3539;
        test_state <= test_b1_S4658;
      end
      test_b1_S4658: begin
        IMAGE_addr <= 4642;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4598;
        test_state <= test_b1_S4659;
      end
      test_b1_S4659: begin
        IMAGE_addr <= 4643;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4533;
        test_state <= test_b1_S4660;
      end
      test_b1_S4660: begin
        IMAGE_addr <= 4644;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4559;
        test_state <= test_b1_S4661;
      end
      test_b1_S4661: begin
        IMAGE_addr <= 4645;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S4662;
      end
      test_b1_S4662: begin
        IMAGE_addr <= 4646;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4473;
        test_state <= test_b1_S4663;
      end
      test_b1_S4663: begin
        IMAGE_addr <= 4647;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4664;
      end
      test_b1_S4664: begin
        IMAGE_addr <= 4648;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4665;
      end
      test_b1_S4665: begin
        IMAGE_addr <= 4649;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4613;
        test_state <= test_b1_S4666;
      end
      test_b1_S4666: begin
        IMAGE_addr <= 4650;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S4667;
      end
      test_b1_S4667: begin
        IMAGE_addr <= 4651;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4658;
        test_state <= test_b1_S4668;
      end
      test_b1_S4668: begin
        IMAGE_addr <= 4652;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 99;
        test_state <= test_b1_S4669;
      end
      test_b1_S4669: begin
        IMAGE_addr <= 4653;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 108;
        test_state <= test_b1_S4670;
      end
      test_b1_S4670: begin
        IMAGE_addr <= 4654;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S4671;
      end
      test_b1_S4671: begin
        IMAGE_addr <= 4655;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S4672;
      end
      test_b1_S4672: begin
        IMAGE_addr <= 4656;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S4673;
      end
      test_b1_S4673: begin
        IMAGE_addr <= 4657;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4674;
      end
      test_b1_S4674: begin
        IMAGE_addr <= 4658;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4675;
      end
      test_b1_S4675: begin
        IMAGE_addr <= 4659;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4676;
      end
      test_b1_S4676: begin
        IMAGE_addr <= 4660;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S4677;
      end
      test_b1_S4677: begin
        IMAGE_addr <= 4661;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4294967295;
        test_state <= test_b1_S4678;
      end
      test_b1_S4678: begin
        IMAGE_addr <= 4662;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 359;
        test_state <= test_b1_S4679;
      end
      test_b1_S4679: begin
        IMAGE_addr <= 4663;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4680;
      end
      test_b1_S4680: begin
        IMAGE_addr <= 4664;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4681;
      end
      test_b1_S4681: begin
        IMAGE_addr <= 4665;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4649;
        test_state <= test_b1_S4682;
      end
      test_b1_S4682: begin
        IMAGE_addr <= 4666;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S4683;
      end
      test_b1_S4683: begin
        IMAGE_addr <= 4667;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4674;
        test_state <= test_b1_S4684;
      end
      test_b1_S4684: begin
        IMAGE_addr <= 4668;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S4685;
      end
      test_b1_S4685: begin
        IMAGE_addr <= 4669;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 112;
        test_state <= test_b1_S4686;
      end
      test_b1_S4686: begin
        IMAGE_addr <= 4670;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S4687;
      end
      test_b1_S4687: begin
        IMAGE_addr <= 4671;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 99;
        test_state <= test_b1_S4688;
      end
      test_b1_S4688: begin
        IMAGE_addr <= 4672;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S4689;
      end
      test_b1_S4689: begin
        IMAGE_addr <= 4673;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4690;
      end
      test_b1_S4690: begin
        IMAGE_addr <= 4674;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4691;
      end
      test_b1_S4691: begin
        IMAGE_addr <= 4675;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4692;
      end
      test_b1_S4692: begin
        IMAGE_addr <= 4676;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S4693;
      end
      test_b1_S4693: begin
        IMAGE_addr <= 4677;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 32;
        test_state <= test_b1_S4694;
      end
      test_b1_S4694: begin
        IMAGE_addr <= 4678;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 359;
        test_state <= test_b1_S4695;
      end
      test_b1_S4695: begin
        IMAGE_addr <= 4679;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4696;
      end
      test_b1_S4696: begin
        IMAGE_addr <= 4680;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4697;
      end
      test_b1_S4697: begin
        IMAGE_addr <= 4681;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4665;
        test_state <= test_b1_S4698;
      end
      test_b1_S4698: begin
        IMAGE_addr <= 4682;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S4699;
      end
      test_b1_S4699: begin
        IMAGE_addr <= 4683;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4689;
        test_state <= test_b1_S4700;
      end
      test_b1_S4700: begin
        IMAGE_addr <= 4684;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 112;
        test_state <= test_b1_S4701;
      end
      test_b1_S4701: begin
        IMAGE_addr <= 4685;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 117;
        test_state <= test_b1_S4702;
      end
      test_b1_S4702: begin
        IMAGE_addr <= 4686;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S4703;
      end
      test_b1_S4703: begin
        IMAGE_addr <= 4687;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 110;
        test_state <= test_b1_S4704;
      end
      test_b1_S4704: begin
        IMAGE_addr <= 4688;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4705;
      end
      test_b1_S4705: begin
        IMAGE_addr <= 4689;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4706;
      end
      test_b1_S4706: begin
        IMAGE_addr <= 4690;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4707;
      end
      test_b1_S4707: begin
        IMAGE_addr <= 4691;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4625;
        test_state <= test_b1_S4708;
      end
      test_b1_S4708: begin
        IMAGE_addr <= 4692;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 391;
        test_state <= test_b1_S4709;
      end
      test_b1_S4709: begin
        IMAGE_addr <= 4693;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4710;
      end
      test_b1_S4710: begin
        IMAGE_addr <= 4694;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4711;
      end
      test_b1_S4711: begin
        IMAGE_addr <= 4695;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4681;
        test_state <= test_b1_S4712;
      end
      test_b1_S4712: begin
        IMAGE_addr <= 4696;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S4713;
      end
      test_b1_S4713: begin
        IMAGE_addr <= 4697;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4705;
        test_state <= test_b1_S4714;
      end
      test_b1_S4714: begin
        IMAGE_addr <= 4698;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 46;
        test_state <= test_b1_S4715;
      end
      test_b1_S4715: begin
        IMAGE_addr <= 4699;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 112;
        test_state <= test_b1_S4716;
      end
      test_b1_S4716: begin
        IMAGE_addr <= 4700;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S4717;
      end
      test_b1_S4717: begin
        IMAGE_addr <= 4701;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S4718;
      end
      test_b1_S4718: begin
        IMAGE_addr <= 4702;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S4719;
      end
      test_b1_S4719: begin
        IMAGE_addr <= 4703;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S4720;
      end
      test_b1_S4720: begin
        IMAGE_addr <= 4704;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4721;
      end
      test_b1_S4721: begin
        IMAGE_addr <= 4705;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4722;
      end
      test_b1_S4722: begin
        IMAGE_addr <= 4706;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4723;
      end
      test_b1_S4723: begin
        IMAGE_addr <= 4707;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 183;
        test_state <= test_b1_S4724;
      end
      test_b1_S4724: begin
        IMAGE_addr <= 4708;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4725;
      end
      test_b1_S4725: begin
        IMAGE_addr <= 4709;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4726;
      end
      test_b1_S4726: begin
        IMAGE_addr <= 4710;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4695;
        test_state <= test_b1_S4727;
      end
      test_b1_S4727: begin
        IMAGE_addr <= 4711;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S4728;
      end
      test_b1_S4728: begin
        IMAGE_addr <= 4712;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4721;
        test_state <= test_b1_S4729;
      end
      test_b1_S4729: begin
        IMAGE_addr <= 4713;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 112;
        test_state <= test_b1_S4730;
      end
      test_b1_S4730: begin
        IMAGE_addr <= 4714;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S4731;
      end
      test_b1_S4731: begin
        IMAGE_addr <= 4715;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S4732;
      end
      test_b1_S4732: begin
        IMAGE_addr <= 4716;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S4733;
      end
      test_b1_S4733: begin
        IMAGE_addr <= 4717;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S4734;
      end
      test_b1_S4734: begin
        IMAGE_addr <= 4718;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 110;
        test_state <= test_b1_S4735;
      end
      test_b1_S4735: begin
        IMAGE_addr <= 4719;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 103;
        test_state <= test_b1_S4736;
      end
      test_b1_S4736: begin
        IMAGE_addr <= 4720;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4737;
      end
      test_b1_S4737: begin
        IMAGE_addr <= 4721;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4738;
      end
      test_b1_S4738: begin
        IMAGE_addr <= 4722;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4739;
      end
      test_b1_S4739: begin
        IMAGE_addr <= 4723;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S4740;
      end
      test_b1_S4740: begin
        IMAGE_addr <= 4724;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4705;
        test_state <= test_b1_S4741;
      end
      test_b1_S4741: begin
        IMAGE_addr <= 4725;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3135;
        test_state <= test_b1_S4742;
      end
      test_b1_S4742: begin
        IMAGE_addr <= 4726;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4743;
      end
      test_b1_S4743: begin
        IMAGE_addr <= 4727;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4744;
      end
      test_b1_S4744: begin
        IMAGE_addr <= 4728;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4710;
        test_state <= test_b1_S4745;
      end
      test_b1_S4745: begin
        IMAGE_addr <= 4729;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S4746;
      end
      test_b1_S4746: begin
        IMAGE_addr <= 4730;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4738;
        test_state <= test_b1_S4747;
      end
      test_b1_S4747: begin
        IMAGE_addr <= 4731;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 110;
        test_state <= test_b1_S4748;
      end
      test_b1_S4748: begin
        IMAGE_addr <= 4732;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 117;
        test_state <= test_b1_S4749;
      end
      test_b1_S4749: begin
        IMAGE_addr <= 4733;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 109;
        test_state <= test_b1_S4750;
      end
      test_b1_S4750: begin
        IMAGE_addr <= 4734;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 98;
        test_state <= test_b1_S4751;
      end
      test_b1_S4751: begin
        IMAGE_addr <= 4735;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S4752;
      end
      test_b1_S4752: begin
        IMAGE_addr <= 4736;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S4753;
      end
      test_b1_S4753: begin
        IMAGE_addr <= 4737;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4754;
      end
      test_b1_S4754: begin
        IMAGE_addr <= 4738;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S4755;
      end
      test_b1_S4755: begin
        IMAGE_addr <= 4739;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 925;
        test_state <= test_b1_S4756;
      end
      test_b1_S4756: begin
        IMAGE_addr <= 4740;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S4757;
      end
      test_b1_S4757: begin
        IMAGE_addr <= 4741;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4746;
        test_state <= test_b1_S4758;
      end
      test_b1_S4758: begin
        IMAGE_addr <= 4742;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 183;
        test_state <= test_b1_S4759;
      end
      test_b1_S4759: begin
        IMAGE_addr <= 4743;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1056;
        test_state <= test_b1_S4760;
      end
      test_b1_S4760: begin
        IMAGE_addr <= 4744;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 310;
        test_state <= test_b1_S4761;
      end
      test_b1_S4761: begin
        IMAGE_addr <= 4745;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4762;
      end
      test_b1_S4762: begin
        IMAGE_addr <= 4746;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3673;
        test_state <= test_b1_S4763;
      end
      test_b1_S4763: begin
        IMAGE_addr <= 4747;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4764;
      end
      test_b1_S4764: begin
        IMAGE_addr <= 4748;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4765;
      end
      test_b1_S4765: begin
        IMAGE_addr <= 4749;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4710;
        test_state <= test_b1_S4766;
      end
      test_b1_S4766: begin
        IMAGE_addr <= 4750;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4705;
        test_state <= test_b1_S4767;
      end
      test_b1_S4767: begin
        IMAGE_addr <= 4751;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4756;
        test_state <= test_b1_S4768;
      end
      test_b1_S4768: begin
        IMAGE_addr <= 4752;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 95;
        test_state <= test_b1_S4769;
      end
      test_b1_S4769: begin
        IMAGE_addr <= 4753;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 95;
        test_state <= test_b1_S4770;
      end
      test_b1_S4770: begin
        IMAGE_addr <= 4754;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 36;
        test_state <= test_b1_S4771;
      end
      test_b1_S4771: begin
        IMAGE_addr <= 4755;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4772;
      end
      test_b1_S4772: begin
        IMAGE_addr <= 4756;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4773;
      end
      test_b1_S4773: begin
        IMAGE_addr <= 4757;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4774;
      end
      test_b1_S4774: begin
        IMAGE_addr <= 4758;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S4775;
      end
      test_b1_S4775: begin
        IMAGE_addr <= 4759;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4420;
        test_state <= test_b1_S4776;
      end
      test_b1_S4776: begin
        IMAGE_addr <= 4760;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4738;
        test_state <= test_b1_S4777;
      end
      test_b1_S4777: begin
        IMAGE_addr <= 4761;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4778;
      end
      test_b1_S4778: begin
        IMAGE_addr <= 4762;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4779;
      end
      test_b1_S4779: begin
        IMAGE_addr <= 4763;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4749;
        test_state <= test_b1_S4780;
      end
      test_b1_S4780: begin
        IMAGE_addr <= 4764;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4705;
        test_state <= test_b1_S4781;
      end
      test_b1_S4781: begin
        IMAGE_addr <= 4765;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4770;
        test_state <= test_b1_S4782;
      end
      test_b1_S4782: begin
        IMAGE_addr <= 4766;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 95;
        test_state <= test_b1_S4783;
      end
      test_b1_S4783: begin
        IMAGE_addr <= 4767;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 95;
        test_state <= test_b1_S4784;
      end
      test_b1_S4784: begin
        IMAGE_addr <= 4768;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 35;
        test_state <= test_b1_S4785;
      end
      test_b1_S4785: begin
        IMAGE_addr <= 4769;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4786;
      end
      test_b1_S4786: begin
        IMAGE_addr <= 4770;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4787;
      end
      test_b1_S4787: begin
        IMAGE_addr <= 4771;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4788;
      end
      test_b1_S4788: begin
        IMAGE_addr <= 4772;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S4789;
      end
      test_b1_S4789: begin
        IMAGE_addr <= 4773;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4404;
        test_state <= test_b1_S4790;
      end
      test_b1_S4790: begin
        IMAGE_addr <= 4774;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4738;
        test_state <= test_b1_S4791;
      end
      test_b1_S4791: begin
        IMAGE_addr <= 4775;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4792;
      end
      test_b1_S4792: begin
        IMAGE_addr <= 4776;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4793;
      end
      test_b1_S4793: begin
        IMAGE_addr <= 4777;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4763;
        test_state <= test_b1_S4794;
      end
      test_b1_S4794: begin
        IMAGE_addr <= 4778;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4705;
        test_state <= test_b1_S4795;
      end
      test_b1_S4795: begin
        IMAGE_addr <= 4779;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4784;
        test_state <= test_b1_S4796;
      end
      test_b1_S4796: begin
        IMAGE_addr <= 4780;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 95;
        test_state <= test_b1_S4797;
      end
      test_b1_S4797: begin
        IMAGE_addr <= 4781;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 95;
        test_state <= test_b1_S4798;
      end
      test_b1_S4798: begin
        IMAGE_addr <= 4782;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 37;
        test_state <= test_b1_S4799;
      end
      test_b1_S4799: begin
        IMAGE_addr <= 4783;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4800;
      end
      test_b1_S4800: begin
        IMAGE_addr <= 4784;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4801;
      end
      test_b1_S4801: begin
        IMAGE_addr <= 4785;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4802;
      end
      test_b1_S4802: begin
        IMAGE_addr <= 4786;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S4803;
      end
      test_b1_S4803: begin
        IMAGE_addr <= 4787;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4457;
        test_state <= test_b1_S4804;
      end
      test_b1_S4804: begin
        IMAGE_addr <= 4788;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4738;
        test_state <= test_b1_S4805;
      end
      test_b1_S4805: begin
        IMAGE_addr <= 4789;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4806;
      end
      test_b1_S4806: begin
        IMAGE_addr <= 4790;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4807;
      end
      test_b1_S4807: begin
        IMAGE_addr <= 4791;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4777;
        test_state <= test_b1_S4808;
      end
      test_b1_S4808: begin
        IMAGE_addr <= 4792;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4705;
        test_state <= test_b1_S4809;
      end
      test_b1_S4809: begin
        IMAGE_addr <= 4793;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4798;
        test_state <= test_b1_S4810;
      end
      test_b1_S4810: begin
        IMAGE_addr <= 4794;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 95;
        test_state <= test_b1_S4811;
      end
      test_b1_S4811: begin
        IMAGE_addr <= 4795;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 95;
        test_state <= test_b1_S4812;
      end
      test_b1_S4812: begin
        IMAGE_addr <= 4796;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 39;
        test_state <= test_b1_S4813;
      end
      test_b1_S4813: begin
        IMAGE_addr <= 4797;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4814;
      end
      test_b1_S4814: begin
        IMAGE_addr <= 4798;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4815;
      end
      test_b1_S4815: begin
        IMAGE_addr <= 4799;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4816;
      end
      test_b1_S4816: begin
        IMAGE_addr <= 4800;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S4817;
      end
      test_b1_S4817: begin
        IMAGE_addr <= 4801;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 310;
        test_state <= test_b1_S4818;
      end
      test_b1_S4818: begin
        IMAGE_addr <= 4802;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4819;
      end
      test_b1_S4819: begin
        IMAGE_addr <= 4803;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4820;
      end
      test_b1_S4820: begin
        IMAGE_addr <= 4804;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4791;
        test_state <= test_b1_S4821;
      end
      test_b1_S4821: begin
        IMAGE_addr <= 4805;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 310;
        test_state <= test_b1_S4822;
      end
      test_b1_S4822: begin
        IMAGE_addr <= 4806;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4813;
        test_state <= test_b1_S4823;
      end
      test_b1_S4823: begin
        IMAGE_addr <= 4807;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 100;
        test_state <= test_b1_S4824;
      end
      test_b1_S4824: begin
        IMAGE_addr <= 4808;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S4825;
      end
      test_b1_S4825: begin
        IMAGE_addr <= 4809;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 99;
        test_state <= test_b1_S4826;
      end
      test_b1_S4826: begin
        IMAGE_addr <= 4810;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S4827;
      end
      test_b1_S4827: begin
        IMAGE_addr <= 4811;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S4828;
      end
      test_b1_S4828: begin
        IMAGE_addr <= 4812;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4829;
      end
      test_b1_S4829: begin
        IMAGE_addr <= 4813;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4830;
      end
      test_b1_S4830: begin
        IMAGE_addr <= 4814;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7933;
        test_state <= test_b1_S4831;
      end
      test_b1_S4831: begin
        IMAGE_addr <= 4815;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4832;
      end
      test_b1_S4832: begin
        IMAGE_addr <= 4816;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4833;
      end
      test_b1_S4833: begin
        IMAGE_addr <= 4817;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4834;
      end
      test_b1_S4834: begin
        IMAGE_addr <= 4818;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4835;
      end
      test_b1_S4835: begin
        IMAGE_addr <= 4819;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4836;
      end
      test_b1_S4836: begin
        IMAGE_addr <= 4820;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4837;
      end
      test_b1_S4837: begin
        IMAGE_addr <= 4821;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4838;
      end
      test_b1_S4838: begin
        IMAGE_addr <= 4822;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4839;
      end
      test_b1_S4839: begin
        IMAGE_addr <= 4823;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4840;
      end
      test_b1_S4840: begin
        IMAGE_addr <= 4824;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4841;
      end
      test_b1_S4841: begin
        IMAGE_addr <= 4825;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4842;
      end
      test_b1_S4842: begin
        IMAGE_addr <= 4826;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4843;
      end
      test_b1_S4843: begin
        IMAGE_addr <= 4827;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4844;
      end
      test_b1_S4844: begin
        IMAGE_addr <= 4828;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4845;
      end
      test_b1_S4845: begin
        IMAGE_addr <= 4829;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4846;
      end
      test_b1_S4846: begin
        IMAGE_addr <= 4830;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4847;
      end
      test_b1_S4847: begin
        IMAGE_addr <= 4831;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4848;
      end
      test_b1_S4848: begin
        IMAGE_addr <= 4832;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4849;
      end
      test_b1_S4849: begin
        IMAGE_addr <= 4833;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4850;
      end
      test_b1_S4850: begin
        IMAGE_addr <= 4834;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4851;
      end
      test_b1_S4851: begin
        IMAGE_addr <= 4835;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4852;
      end
      test_b1_S4852: begin
        IMAGE_addr <= 4836;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4853;
      end
      test_b1_S4853: begin
        IMAGE_addr <= 4837;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4854;
      end
      test_b1_S4854: begin
        IMAGE_addr <= 4838;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4855;
      end
      test_b1_S4855: begin
        IMAGE_addr <= 4839;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4856;
      end
      test_b1_S4856: begin
        IMAGE_addr <= 4840;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4857;
      end
      test_b1_S4857: begin
        IMAGE_addr <= 4841;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4858;
      end
      test_b1_S4858: begin
        IMAGE_addr <= 4842;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4859;
      end
      test_b1_S4859: begin
        IMAGE_addr <= 4843;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4860;
      end
      test_b1_S4860: begin
        IMAGE_addr <= 4844;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4861;
      end
      test_b1_S4861: begin
        IMAGE_addr <= 4845;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4862;
      end
      test_b1_S4862: begin
        IMAGE_addr <= 4846;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4863;
      end
      test_b1_S4863: begin
        IMAGE_addr <= 4847;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4864;
      end
      test_b1_S4864: begin
        IMAGE_addr <= 4848;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4865;
      end
      test_b1_S4865: begin
        IMAGE_addr <= 4849;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4866;
      end
      test_b1_S4866: begin
        IMAGE_addr <= 4850;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4867;
      end
      test_b1_S4867: begin
        IMAGE_addr <= 4851;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4868;
      end
      test_b1_S4868: begin
        IMAGE_addr <= 4852;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4869;
      end
      test_b1_S4869: begin
        IMAGE_addr <= 4853;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4870;
      end
      test_b1_S4870: begin
        IMAGE_addr <= 4854;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4871;
      end
      test_b1_S4871: begin
        IMAGE_addr <= 4855;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4872;
      end
      test_b1_S4872: begin
        IMAGE_addr <= 4856;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4873;
      end
      test_b1_S4873: begin
        IMAGE_addr <= 4857;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4874;
      end
      test_b1_S4874: begin
        IMAGE_addr <= 4858;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4875;
      end
      test_b1_S4875: begin
        IMAGE_addr <= 4859;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4876;
      end
      test_b1_S4876: begin
        IMAGE_addr <= 4860;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4877;
      end
      test_b1_S4877: begin
        IMAGE_addr <= 4861;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4878;
      end
      test_b1_S4878: begin
        IMAGE_addr <= 4862;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4879;
      end
      test_b1_S4879: begin
        IMAGE_addr <= 4863;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4880;
      end
      test_b1_S4880: begin
        IMAGE_addr <= 4864;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4881;
      end
      test_b1_S4881: begin
        IMAGE_addr <= 4865;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4882;
      end
      test_b1_S4882: begin
        IMAGE_addr <= 4866;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4883;
      end
      test_b1_S4883: begin
        IMAGE_addr <= 4867;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4884;
      end
      test_b1_S4884: begin
        IMAGE_addr <= 4868;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4885;
      end
      test_b1_S4885: begin
        IMAGE_addr <= 4869;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4886;
      end
      test_b1_S4886: begin
        IMAGE_addr <= 4870;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4887;
      end
      test_b1_S4887: begin
        IMAGE_addr <= 4871;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4888;
      end
      test_b1_S4888: begin
        IMAGE_addr <= 4872;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4889;
      end
      test_b1_S4889: begin
        IMAGE_addr <= 4873;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4890;
      end
      test_b1_S4890: begin
        IMAGE_addr <= 4874;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4891;
      end
      test_b1_S4891: begin
        IMAGE_addr <= 4875;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4892;
      end
      test_b1_S4892: begin
        IMAGE_addr <= 4876;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4893;
      end
      test_b1_S4893: begin
        IMAGE_addr <= 4877;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8479;
        test_state <= test_b1_S4894;
      end
      test_b1_S4894: begin
        IMAGE_addr <= 4878;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8004;
        test_state <= test_b1_S4895;
      end
      test_b1_S4895: begin
        IMAGE_addr <= 4879;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4804;
        test_state <= test_b1_S4896;
      end
      test_b1_S4896: begin
        IMAGE_addr <= 4880;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 310;
        test_state <= test_b1_S4897;
      end
      test_b1_S4897: begin
        IMAGE_addr <= 4881;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4877;
        test_state <= test_b1_S4898;
      end
      test_b1_S4898: begin
        IMAGE_addr <= 4882;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S4899;
      end
      test_b1_S4899: begin
        IMAGE_addr <= 4883;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 99;
        test_state <= test_b1_S4900;
      end
      test_b1_S4900: begin
        IMAGE_addr <= 4884;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S4901;
      end
      test_b1_S4901: begin
        IMAGE_addr <= 4885;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S4902;
      end
      test_b1_S4902: begin
        IMAGE_addr <= 4886;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 118;
        test_state <= test_b1_S4903;
      end
      test_b1_S4903: begin
        IMAGE_addr <= 4887;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S4904;
      end
      test_b1_S4904: begin
        IMAGE_addr <= 4888;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4905;
      end
      test_b1_S4905: begin
        IMAGE_addr <= 4889;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4879;
        test_state <= test_b1_S4906;
      end
      test_b1_S4906: begin
        IMAGE_addr <= 4890;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 310;
        test_state <= test_b1_S4907;
      end
      test_b1_S4907: begin
        IMAGE_addr <= 4891;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4878;
        test_state <= test_b1_S4908;
      end
      test_b1_S4908: begin
        IMAGE_addr <= 4892;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 112;
        test_state <= test_b1_S4909;
      end
      test_b1_S4909: begin
        IMAGE_addr <= 4893;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S4910;
      end
      test_b1_S4910: begin
        IMAGE_addr <= 4894;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S4911;
      end
      test_b1_S4911: begin
        IMAGE_addr <= 4895;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 111;
        test_state <= test_b1_S4912;
      end
      test_b1_S4912: begin
        IMAGE_addr <= 4896;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S4913;
      end
      test_b1_S4913: begin
        IMAGE_addr <= 4897;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4914;
      end
      test_b1_S4914: begin
        IMAGE_addr <= 4898;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4889;
        test_state <= test_b1_S4915;
      end
      test_b1_S4915: begin
        IMAGE_addr <= 4899;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 310;
        test_state <= test_b1_S4916;
      end
      test_b1_S4916: begin
        IMAGE_addr <= 4900;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4905;
        test_state <= test_b1_S4917;
      end
      test_b1_S4917: begin
        IMAGE_addr <= 4901;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 34;
        test_state <= test_b1_S4918;
      end
      test_b1_S4918: begin
        IMAGE_addr <= 4902;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 124;
        test_state <= test_b1_S4919;
      end
      test_b1_S4919: begin
        IMAGE_addr <= 4903;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 34;
        test_state <= test_b1_S4920;
      end
      test_b1_S4920: begin
        IMAGE_addr <= 4904;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4921;
      end
      test_b1_S4921: begin
        IMAGE_addr <= 4905;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 124;
        test_state <= test_b1_S4922;
      end
      test_b1_S4922: begin
        IMAGE_addr <= 4906;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4923;
      end
      test_b1_S4923: begin
        IMAGE_addr <= 4907;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4898;
        test_state <= test_b1_S4924;
      end
      test_b1_S4924: begin
        IMAGE_addr <= 4908;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 310;
        test_state <= test_b1_S4925;
      end
      test_b1_S4925: begin
        IMAGE_addr <= 4909;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4915;
        test_state <= test_b1_S4926;
      end
      test_b1_S4926: begin
        IMAGE_addr <= 4910;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 34;
        test_state <= test_b1_S4927;
      end
      test_b1_S4927: begin
        IMAGE_addr <= 4911;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 37;
        test_state <= test_b1_S4928;
      end
      test_b1_S4928: begin
        IMAGE_addr <= 4912;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 37;
        test_state <= test_b1_S4929;
      end
      test_b1_S4929: begin
        IMAGE_addr <= 4913;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 34;
        test_state <= test_b1_S4930;
      end
      test_b1_S4930: begin
        IMAGE_addr <= 4914;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4931;
      end
      test_b1_S4931: begin
        IMAGE_addr <= 4915;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 37;
        test_state <= test_b1_S4932;
      end
      test_b1_S4932: begin
        IMAGE_addr <= 4916;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 37;
        test_state <= test_b1_S4933;
      end
      test_b1_S4933: begin
        IMAGE_addr <= 4917;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4934;
      end
      test_b1_S4934: begin
        IMAGE_addr <= 4918;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4907;
        test_state <= test_b1_S4935;
      end
      test_b1_S4935: begin
        IMAGE_addr <= 4919;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S4936;
      end
      test_b1_S4936: begin
        IMAGE_addr <= 4920;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4926;
        test_state <= test_b1_S4937;
      end
      test_b1_S4937: begin
        IMAGE_addr <= 4921;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S4938;
      end
      test_b1_S4938: begin
        IMAGE_addr <= 4922;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S4939;
      end
      test_b1_S4939: begin
        IMAGE_addr <= 4923;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S4940;
      end
      test_b1_S4940: begin
        IMAGE_addr <= 4924;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 108;
        test_state <= test_b1_S4941;
      end
      test_b1_S4941: begin
        IMAGE_addr <= 4925;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4942;
      end
      test_b1_S4942: begin
        IMAGE_addr <= 4926;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S4943;
      end
      test_b1_S4943: begin
        IMAGE_addr <= 4927;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S4944;
      end
      test_b1_S4944: begin
        IMAGE_addr <= 4928;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S4945;
      end
      test_b1_S4945: begin
        IMAGE_addr <= 4929;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4939;
        test_state <= test_b1_S4946;
      end
      test_b1_S4946: begin
        IMAGE_addr <= 4930;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S4947;
      end
      test_b1_S4947: begin
        IMAGE_addr <= 4931;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 25;
        test_state <= test_b1_S4948;
      end
      test_b1_S4948: begin
        IMAGE_addr <= 4932;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S4949;
      end
      test_b1_S4949: begin
        IMAGE_addr <= 4933;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4877;
        test_state <= test_b1_S4950;
      end
      test_b1_S4950: begin
        IMAGE_addr <= 4934;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S4951;
      end
      test_b1_S4951: begin
        IMAGE_addr <= 4935;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 132;
        test_state <= test_b1_S4952;
      end
      test_b1_S4952: begin
        IMAGE_addr <= 4936;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S4953;
      end
      test_b1_S4953: begin
        IMAGE_addr <= 4937;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 790;
        test_state <= test_b1_S4954;
      end
      test_b1_S4954: begin
        IMAGE_addr <= 4938;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4955;
      end
      test_b1_S4955: begin
        IMAGE_addr <= 4939;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3458;
        test_state <= test_b1_S4956;
      end
      test_b1_S4956: begin
        IMAGE_addr <= 4940;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S4957;
      end
      test_b1_S4957: begin
        IMAGE_addr <= 4941;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4958;
      end
      test_b1_S4958: begin
        IMAGE_addr <= 4942;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S4959;
      end
      test_b1_S4959: begin
        IMAGE_addr <= 4943;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S4960;
      end
      test_b1_S4960: begin
        IMAGE_addr <= 4944;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4961;
      end
      test_b1_S4961: begin
        IMAGE_addr <= 4945;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4962;
      end
      test_b1_S4962: begin
        IMAGE_addr <= 4946;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4918;
        test_state <= test_b1_S4963;
      end
      test_b1_S4963: begin
        IMAGE_addr <= 4947;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S4964;
      end
      test_b1_S4964: begin
        IMAGE_addr <= 4948;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4956;
        test_state <= test_b1_S4965;
      end
      test_b1_S4965: begin
        IMAGE_addr <= 4949;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S4966;
      end
      test_b1_S4966: begin
        IMAGE_addr <= 4950;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S4967;
      end
      test_b1_S4967: begin
        IMAGE_addr <= 4951;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 118;
        test_state <= test_b1_S4968;
      end
      test_b1_S4968: begin
        IMAGE_addr <= 4952;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S4969;
      end
      test_b1_S4969: begin
        IMAGE_addr <= 4953;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S4970;
      end
      test_b1_S4970: begin
        IMAGE_addr <= 4954;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S4971;
      end
      test_b1_S4971: begin
        IMAGE_addr <= 4955;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4972;
      end
      test_b1_S4972: begin
        IMAGE_addr <= 4956;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S4973;
      end
      test_b1_S4973: begin
        IMAGE_addr <= 4957;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4878;
        test_state <= test_b1_S4974;
      end
      test_b1_S4974: begin
        IMAGE_addr <= 4958;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S4975;
      end
      test_b1_S4975: begin
        IMAGE_addr <= 4959;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 25;
        test_state <= test_b1_S4976;
      end
      test_b1_S4976: begin
        IMAGE_addr <= 4960;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S4977;
      end
      test_b1_S4977: begin
        IMAGE_addr <= 4961;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S4978;
      end
      test_b1_S4978: begin
        IMAGE_addr <= 4962;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S4979;
      end
      test_b1_S4979: begin
        IMAGE_addr <= 4963;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S4980;
      end
      test_b1_S4980: begin
        IMAGE_addr <= 4964;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4981;
      end
      test_b1_S4981: begin
        IMAGE_addr <= 4965;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S4982;
      end
      test_b1_S4982: begin
        IMAGE_addr <= 4966;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4878;
        test_state <= test_b1_S4983;
      end
      test_b1_S4983: begin
        IMAGE_addr <= 4967;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S4984;
      end
      test_b1_S4984: begin
        IMAGE_addr <= 4968;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4985;
      end
      test_b1_S4985: begin
        IMAGE_addr <= 4969;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S4986;
      end
      test_b1_S4986: begin
        IMAGE_addr <= 4970;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4946;
        test_state <= test_b1_S4987;
      end
      test_b1_S4987: begin
        IMAGE_addr <= 4971;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S4988;
      end
      test_b1_S4988: begin
        IMAGE_addr <= 4972;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4980;
        test_state <= test_b1_S4989;
      end
      test_b1_S4989: begin
        IMAGE_addr <= 4973;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S4990;
      end
      test_b1_S4990: begin
        IMAGE_addr <= 4974;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S4991;
      end
      test_b1_S4991: begin
        IMAGE_addr <= 4975;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 102;
        test_state <= test_b1_S4992;
      end
      test_b1_S4992: begin
        IMAGE_addr <= 4976;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S4993;
      end
      test_b1_S4993: begin
        IMAGE_addr <= 4977;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S4994;
      end
      test_b1_S4994: begin
        IMAGE_addr <= 4978;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 121;
        test_state <= test_b1_S4995;
      end
      test_b1_S4995: begin
        IMAGE_addr <= 4979;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S4996;
      end
      test_b1_S4996: begin
        IMAGE_addr <= 4980;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S4997;
      end
      test_b1_S4997: begin
        IMAGE_addr <= 4981;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4915;
        test_state <= test_b1_S4998;
      end
      test_b1_S4998: begin
        IMAGE_addr <= 4982;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 596;
        test_state <= test_b1_S4999;
      end
      test_b1_S4999: begin
        IMAGE_addr <= 4983;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3308;
        test_state <= test_b1_S5000;
      end
      test_b1_S5000: begin
        IMAGE_addr <= 4984;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5001;
      end
      test_b1_S5001: begin
        IMAGE_addr <= 4985;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4956;
        test_state <= test_b1_S5002;
      end
      test_b1_S5002: begin
        IMAGE_addr <= 4986;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5003;
      end
      test_b1_S5003: begin
        IMAGE_addr <= 4987;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S5004;
      end
      test_b1_S5004: begin
        IMAGE_addr <= 4988;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S5005;
      end
      test_b1_S5005: begin
        IMAGE_addr <= 4989;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 583;
        test_state <= test_b1_S5006;
      end
      test_b1_S5006: begin
        IMAGE_addr <= 4990;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S5007;
      end
      test_b1_S5007: begin
        IMAGE_addr <= 4991;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5008;
      end
      test_b1_S5008: begin
        IMAGE_addr <= 4992;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5009;
      end
      test_b1_S5009: begin
        IMAGE_addr <= 4993;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4804;
        test_state <= test_b1_S5010;
      end
      test_b1_S5010: begin
        IMAGE_addr <= 4994;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S5011;
      end
      test_b1_S5011: begin
        IMAGE_addr <= 4995;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4999;
        test_state <= test_b1_S5012;
      end
      test_b1_S5012: begin
        IMAGE_addr <= 4996;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 37;
        test_state <= test_b1_S5013;
      end
      test_b1_S5013: begin
        IMAGE_addr <= 4997;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 37;
        test_state <= test_b1_S5014;
      end
      test_b1_S5014: begin
        IMAGE_addr <= 4998;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S5015;
      end
      test_b1_S5015: begin
        IMAGE_addr <= 4999;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S5016;
      end
      test_b1_S5016: begin
        IMAGE_addr <= 5000;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S5017;
      end
      test_b1_S5017: begin
        IMAGE_addr <= 5001;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4956;
        test_state <= test_b1_S5018;
      end
      test_b1_S5018: begin
        IMAGE_addr <= 5002;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5019;
      end
      test_b1_S5019: begin
        IMAGE_addr <= 5003;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5020;
      end
      test_b1_S5020: begin
        IMAGE_addr <= 5004;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4993;
        test_state <= test_b1_S5021;
      end
      test_b1_S5021: begin
        IMAGE_addr <= 5005;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S5022;
      end
      test_b1_S5022: begin
        IMAGE_addr <= 5006;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5011;
        test_state <= test_b1_S5023;
      end
      test_b1_S5023: begin
        IMAGE_addr <= 5007;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 60;
        test_state <= test_b1_S5024;
      end
      test_b1_S5024: begin
        IMAGE_addr <= 5008;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 37;
        test_state <= test_b1_S5025;
      end
      test_b1_S5025: begin
        IMAGE_addr <= 5009;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 62;
        test_state <= test_b1_S5026;
      end
      test_b1_S5026: begin
        IMAGE_addr <= 5010;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S5027;
      end
      test_b1_S5027: begin
        IMAGE_addr <= 5011;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S5028;
      end
      test_b1_S5028: begin
        IMAGE_addr <= 5012;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S5029;
      end
      test_b1_S5029: begin
        IMAGE_addr <= 5013;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5030;
      end
      test_b1_S5030: begin
        IMAGE_addr <= 5014;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S5031;
      end
      test_b1_S5031: begin
        IMAGE_addr <= 5015;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S5032;
      end
      test_b1_S5032: begin
        IMAGE_addr <= 5016;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5033;
      end
      test_b1_S5033: begin
        IMAGE_addr <= 5017;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4878;
        test_state <= test_b1_S5034;
      end
      test_b1_S5034: begin
        IMAGE_addr <= 5018;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S5035;
      end
      test_b1_S5035: begin
        IMAGE_addr <= 5019;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5036;
      end
      test_b1_S5036: begin
        IMAGE_addr <= 5020;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S5037;
      end
      test_b1_S5037: begin
        IMAGE_addr <= 5021;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S5038;
      end
      test_b1_S5038: begin
        IMAGE_addr <= 5022;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5039;
      end
      test_b1_S5039: begin
        IMAGE_addr <= 5023;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5040;
      end
      test_b1_S5040: begin
        IMAGE_addr <= 5024;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5004;
        test_state <= test_b1_S5041;
      end
      test_b1_S5041: begin
        IMAGE_addr <= 5025;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S5042;
      end
      test_b1_S5042: begin
        IMAGE_addr <= 5026;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5034;
        test_state <= test_b1_S5043;
      end
      test_b1_S5043: begin
        IMAGE_addr <= 5027;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 46;
        test_state <= test_b1_S5044;
      end
      test_b1_S5044: begin
        IMAGE_addr <= 5028;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 99;
        test_state <= test_b1_S5045;
      end
      test_b1_S5045: begin
        IMAGE_addr <= 5029;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 104;
        test_state <= test_b1_S5046;
      end
      test_b1_S5046: begin
        IMAGE_addr <= 5030;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S5047;
      end
      test_b1_S5047: begin
        IMAGE_addr <= 5031;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S5048;
      end
      test_b1_S5048: begin
        IMAGE_addr <= 5032;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 110;
        test_state <= test_b1_S5049;
      end
      test_b1_S5049: begin
        IMAGE_addr <= 5033;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S5050;
      end
      test_b1_S5050: begin
        IMAGE_addr <= 5034;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S5051;
      end
      test_b1_S5051: begin
        IMAGE_addr <= 5035;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S5052;
      end
      test_b1_S5052: begin
        IMAGE_addr <= 5036;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5053;
      end
      test_b1_S5053: begin
        IMAGE_addr <= 5037;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4813;
        test_state <= test_b1_S5054;
      end
      test_b1_S5054: begin
        IMAGE_addr <= 5038;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S5055;
      end
      test_b1_S5055: begin
        IMAGE_addr <= 5039;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5056;
      end
      test_b1_S5056: begin
        IMAGE_addr <= 5040;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 52;
        test_state <= test_b1_S5057;
      end
      test_b1_S5057: begin
        IMAGE_addr <= 5041;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5058;
      end
      test_b1_S5058: begin
        IMAGE_addr <= 5042;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5011;
        test_state <= test_b1_S5059;
      end
      test_b1_S5059: begin
        IMAGE_addr <= 5043;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 732;
        test_state <= test_b1_S5060;
      end
      test_b1_S5060: begin
        IMAGE_addr <= 5044;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5061;
      end
      test_b1_S5061: begin
        IMAGE_addr <= 5045;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5062;
      end
      test_b1_S5062: begin
        IMAGE_addr <= 5046;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5024;
        test_state <= test_b1_S5063;
      end
      test_b1_S5063: begin
        IMAGE_addr <= 5047;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S5064;
      end
      test_b1_S5064: begin
        IMAGE_addr <= 5048;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5056;
        test_state <= test_b1_S5065;
      end
      test_b1_S5065: begin
        IMAGE_addr <= 5049;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 99;
        test_state <= test_b1_S5066;
      end
      test_b1_S5066: begin
        IMAGE_addr <= 5050;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 104;
        test_state <= test_b1_S5067;
      end
      test_b1_S5067: begin
        IMAGE_addr <= 5051;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S5068;
      end
      test_b1_S5068: begin
        IMAGE_addr <= 5052;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S5069;
      end
      test_b1_S5069: begin
        IMAGE_addr <= 5053;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 110;
        test_state <= test_b1_S5070;
      end
      test_b1_S5070: begin
        IMAGE_addr <= 5054;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 58;
        test_state <= test_b1_S5071;
      end
      test_b1_S5071: begin
        IMAGE_addr <= 5055;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S5072;
      end
      test_b1_S5072: begin
        IMAGE_addr <= 5056;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S5073;
      end
      test_b1_S5073: begin
        IMAGE_addr <= 5057;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S5074;
      end
      test_b1_S5074: begin
        IMAGE_addr <= 5058;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 621;
        test_state <= test_b1_S5075;
      end
      test_b1_S5075: begin
        IMAGE_addr <= 5059;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5076;
      end
      test_b1_S5076: begin
        IMAGE_addr <= 5060;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S5077;
      end
      test_b1_S5077: begin
        IMAGE_addr <= 5061;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 213;
        test_state <= test_b1_S5078;
      end
      test_b1_S5078: begin
        IMAGE_addr <= 5062;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5079;
      end
      test_b1_S5079: begin
        IMAGE_addr <= 5063;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5034;
        test_state <= test_b1_S5080;
      end
      test_b1_S5080: begin
        IMAGE_addr <= 5064;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3135;
        test_state <= test_b1_S5081;
      end
      test_b1_S5081: begin
        IMAGE_addr <= 5065;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5082;
      end
      test_b1_S5082: begin
        IMAGE_addr <= 5066;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S5083;
      end
      test_b1_S5083: begin
        IMAGE_addr <= 5067;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S5084;
      end
      test_b1_S5084: begin
        IMAGE_addr <= 5068;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5085;
      end
      test_b1_S5085: begin
        IMAGE_addr <= 5069;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4877;
        test_state <= test_b1_S5086;
      end
      test_b1_S5086: begin
        IMAGE_addr <= 5070;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S5087;
      end
      test_b1_S5087: begin
        IMAGE_addr <= 5071;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4980;
        test_state <= test_b1_S5088;
      end
      test_b1_S5088: begin
        IMAGE_addr <= 5072;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5089;
      end
      test_b1_S5089: begin
        IMAGE_addr <= 5073;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5090;
      end
      test_b1_S5090: begin
        IMAGE_addr <= 5074;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5046;
        test_state <= test_b1_S5091;
      end
      test_b1_S5091: begin
        IMAGE_addr <= 5075;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S5092;
      end
      test_b1_S5092: begin
        IMAGE_addr <= 5076;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5084;
        test_state <= test_b1_S5093;
      end
      test_b1_S5093: begin
        IMAGE_addr <= 5077;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 59;
        test_state <= test_b1_S5094;
      end
      test_b1_S5094: begin
        IMAGE_addr <= 5078;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 99;
        test_state <= test_b1_S5095;
      end
      test_b1_S5095: begin
        IMAGE_addr <= 5079;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 104;
        test_state <= test_b1_S5096;
      end
      test_b1_S5096: begin
        IMAGE_addr <= 5080;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S5097;
      end
      test_b1_S5097: begin
        IMAGE_addr <= 5081;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S5098;
      end
      test_b1_S5098: begin
        IMAGE_addr <= 5082;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 110;
        test_state <= test_b1_S5099;
      end
      test_b1_S5099: begin
        IMAGE_addr <= 5083;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S5100;
      end
      test_b1_S5100: begin
        IMAGE_addr <= 5084;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S5101;
      end
      test_b1_S5101: begin
        IMAGE_addr <= 5085;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S5102;
      end
      test_b1_S5102: begin
        IMAGE_addr <= 5086;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4926;
        test_state <= test_b1_S5103;
      end
      test_b1_S5103: begin
        IMAGE_addr <= 5087;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5104;
      end
      test_b1_S5104: begin
        IMAGE_addr <= 5088;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S5105;
      end
      test_b1_S5105: begin
        IMAGE_addr <= 5089;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S5106;
      end
      test_b1_S5106: begin
        IMAGE_addr <= 5090;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5107;
      end
      test_b1_S5107: begin
        IMAGE_addr <= 5091;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4877;
        test_state <= test_b1_S5108;
      end
      test_b1_S5108: begin
        IMAGE_addr <= 5092;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S5109;
      end
      test_b1_S5109: begin
        IMAGE_addr <= 5093;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S5110;
      end
      test_b1_S5110: begin
        IMAGE_addr <= 5094;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5099;
        test_state <= test_b1_S5111;
      end
      test_b1_S5111: begin
        IMAGE_addr <= 5095;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5112;
      end
      test_b1_S5112: begin
        IMAGE_addr <= 5096;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S5113;
      end
      test_b1_S5113: begin
        IMAGE_addr <= 5097;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S5114;
      end
      test_b1_S5114: begin
        IMAGE_addr <= 5098;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5115;
      end
      test_b1_S5115: begin
        IMAGE_addr <= 5099;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S5116;
      end
      test_b1_S5116: begin
        IMAGE_addr <= 5100;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5104;
        test_state <= test_b1_S5117;
      end
      test_b1_S5117: begin
        IMAGE_addr <= 5101;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 583;
        test_state <= test_b1_S5118;
      end
      test_b1_S5118: begin
        IMAGE_addr <= 5102;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S5119;
      end
      test_b1_S5119: begin
        IMAGE_addr <= 5103;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5120;
      end
      test_b1_S5120: begin
        IMAGE_addr <= 5104;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3539;
        test_state <= test_b1_S5121;
      end
      test_b1_S5121: begin
        IMAGE_addr <= 5105;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5122;
      end
      test_b1_S5122: begin
        IMAGE_addr <= 5106;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5123;
      end
      test_b1_S5123: begin
        IMAGE_addr <= 5107;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5074;
        test_state <= test_b1_S5124;
      end
      test_b1_S5124: begin
        IMAGE_addr <= 5108;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S5125;
      end
      test_b1_S5125: begin
        IMAGE_addr <= 5109;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5116;
        test_state <= test_b1_S5126;
      end
      test_b1_S5126: begin
        IMAGE_addr <= 5110;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 58;
        test_state <= test_b1_S5127;
      end
      test_b1_S5127: begin
        IMAGE_addr <= 5111;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 119;
        test_state <= test_b1_S5128;
      end
      test_b1_S5128: begin
        IMAGE_addr <= 5112;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S5129;
      end
      test_b1_S5129: begin
        IMAGE_addr <= 5113;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S5130;
      end
      test_b1_S5130: begin
        IMAGE_addr <= 5114;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 104;
        test_state <= test_b1_S5131;
      end
      test_b1_S5131: begin
        IMAGE_addr <= 5115;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S5132;
      end
      test_b1_S5132: begin
        IMAGE_addr <= 5116;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S5133;
      end
      test_b1_S5133: begin
        IMAGE_addr <= 5117;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S5134;
      end
      test_b1_S5134: begin
        IMAGE_addr <= 5118;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 25;
        test_state <= test_b1_S5135;
      end
      test_b1_S5135: begin
        IMAGE_addr <= 5119;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5136;
      end
      test_b1_S5136: begin
        IMAGE_addr <= 5120;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4813;
        test_state <= test_b1_S5137;
      end
      test_b1_S5137: begin
        IMAGE_addr <= 5121;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S5138;
      end
      test_b1_S5138: begin
        IMAGE_addr <= 5122;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 26;
        test_state <= test_b1_S5139;
      end
      test_b1_S5139: begin
        IMAGE_addr <= 5123;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5140;
      end
      test_b1_S5140: begin
        IMAGE_addr <= 5124;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4813;
        test_state <= test_b1_S5141;
      end
      test_b1_S5141: begin
        IMAGE_addr <= 5125;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 16;
        test_state <= test_b1_S5142;
      end
      test_b1_S5142: begin
        IMAGE_addr <= 5126;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S5143;
      end
      test_b1_S5143: begin
        IMAGE_addr <= 5127;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5144;
      end
      test_b1_S5144: begin
        IMAGE_addr <= 5128;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4813;
        test_state <= test_b1_S5145;
      end
      test_b1_S5145: begin
        IMAGE_addr <= 5129;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2651;
        test_state <= test_b1_S5146;
      end
      test_b1_S5146: begin
        IMAGE_addr <= 5130;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5147;
      end
      test_b1_S5147: begin
        IMAGE_addr <= 5131;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5148;
      end
      test_b1_S5148: begin
        IMAGE_addr <= 5132;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5107;
        test_state <= test_b1_S5149;
      end
      test_b1_S5149: begin
        IMAGE_addr <= 5133;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S5150;
      end
      test_b1_S5150: begin
        IMAGE_addr <= 5134;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5140;
        test_state <= test_b1_S5151;
      end
      test_b1_S5151: begin
        IMAGE_addr <= 5135;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 119;
        test_state <= test_b1_S5152;
      end
      test_b1_S5152: begin
        IMAGE_addr <= 5136;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S5153;
      end
      test_b1_S5153: begin
        IMAGE_addr <= 5137;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S5154;
      end
      test_b1_S5154: begin
        IMAGE_addr <= 5138;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 104;
        test_state <= test_b1_S5155;
      end
      test_b1_S5155: begin
        IMAGE_addr <= 5139;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S5156;
      end
      test_b1_S5156: begin
        IMAGE_addr <= 5140;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S5157;
      end
      test_b1_S5157: begin
        IMAGE_addr <= 5141;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S5158;
      end
      test_b1_S5158: begin
        IMAGE_addr <= 5142;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1239;
        test_state <= test_b1_S5159;
      end
      test_b1_S5159: begin
        IMAGE_addr <= 5143;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5116;
        test_state <= test_b1_S5160;
      end
      test_b1_S5160: begin
        IMAGE_addr <= 5144;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5161;
      end
      test_b1_S5161: begin
        IMAGE_addr <= 5145;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5162;
      end
      test_b1_S5162: begin
        IMAGE_addr <= 5146;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5132;
        test_state <= test_b1_S5163;
      end
      test_b1_S5163: begin
        IMAGE_addr <= 5147;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S5164;
      end
      test_b1_S5164: begin
        IMAGE_addr <= 5148;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5157;
        test_state <= test_b1_S5165;
      end
      test_b1_S5165: begin
        IMAGE_addr <= 5149;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 119;
        test_state <= test_b1_S5166;
      end
      test_b1_S5166: begin
        IMAGE_addr <= 5150;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S5167;
      end
      test_b1_S5167: begin
        IMAGE_addr <= 5151;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S5168;
      end
      test_b1_S5168: begin
        IMAGE_addr <= 5152;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 104;
        test_state <= test_b1_S5169;
      end
      test_b1_S5169: begin
        IMAGE_addr <= 5153;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 111;
        test_state <= test_b1_S5170;
      end
      test_b1_S5170: begin
        IMAGE_addr <= 5154;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 117;
        test_state <= test_b1_S5171;
      end
      test_b1_S5171: begin
        IMAGE_addr <= 5155;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S5172;
      end
      test_b1_S5172: begin
        IMAGE_addr <= 5156;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S5173;
      end
      test_b1_S5173: begin
        IMAGE_addr <= 5157;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S5174;
      end
      test_b1_S5174: begin
        IMAGE_addr <= 5158;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S5175;
      end
      test_b1_S5175: begin
        IMAGE_addr <= 5159;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5176;
      end
      test_b1_S5176: begin
        IMAGE_addr <= 5160;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4813;
        test_state <= test_b1_S5177;
      end
      test_b1_S5177: begin
        IMAGE_addr <= 5161;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S5178;
      end
      test_b1_S5178: begin
        IMAGE_addr <= 5162;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 25;
        test_state <= test_b1_S5179;
      end
      test_b1_S5179: begin
        IMAGE_addr <= 5163;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 27;
        test_state <= test_b1_S5180;
      end
      test_b1_S5180: begin
        IMAGE_addr <= 5164;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5181;
      end
      test_b1_S5181: begin
        IMAGE_addr <= 5165;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4813;
        test_state <= test_b1_S5182;
      end
      test_b1_S5182: begin
        IMAGE_addr <= 5166;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S5183;
      end
      test_b1_S5183: begin
        IMAGE_addr <= 5167;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5184;
      end
      test_b1_S5184: begin
        IMAGE_addr <= 5168;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5185;
      end
      test_b1_S5185: begin
        IMAGE_addr <= 5169;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5146;
        test_state <= test_b1_S5186;
      end
      test_b1_S5186: begin
        IMAGE_addr <= 5170;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S5187;
      end
      test_b1_S5187: begin
        IMAGE_addr <= 5171;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5179;
        test_state <= test_b1_S5188;
      end
      test_b1_S5188: begin
        IMAGE_addr <= 5172;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 103;
        test_state <= test_b1_S5189;
      end
      test_b1_S5189: begin
        IMAGE_addr <= 5173;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 108;
        test_state <= test_b1_S5190;
      end
      test_b1_S5190: begin
        IMAGE_addr <= 5174;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 111;
        test_state <= test_b1_S5191;
      end
      test_b1_S5191: begin
        IMAGE_addr <= 5175;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 98;
        test_state <= test_b1_S5192;
      end
      test_b1_S5192: begin
        IMAGE_addr <= 5176;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S5193;
      end
      test_b1_S5193: begin
        IMAGE_addr <= 5177;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 108;
        test_state <= test_b1_S5194;
      end
      test_b1_S5194: begin
        IMAGE_addr <= 5178;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S5195;
      end
      test_b1_S5195: begin
        IMAGE_addr <= 5179;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S5196;
      end
      test_b1_S5196: begin
        IMAGE_addr <= 5180;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S5197;
      end
      test_b1_S5197: begin
        IMAGE_addr <= 5181;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5198;
      end
      test_b1_S5198: begin
        IMAGE_addr <= 5182;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S5199;
      end
      test_b1_S5199: begin
        IMAGE_addr <= 5183;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5200;
      end
      test_b1_S5200: begin
        IMAGE_addr <= 5184;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4813;
        test_state <= test_b1_S5201;
      end
      test_b1_S5201: begin
        IMAGE_addr <= 5185;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S5202;
      end
      test_b1_S5202: begin
        IMAGE_addr <= 5186;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5203;
      end
      test_b1_S5203: begin
        IMAGE_addr <= 5187;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5204;
      end
      test_b1_S5204: begin
        IMAGE_addr <= 5188;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5169;
        test_state <= test_b1_S5205;
      end
      test_b1_S5205: begin
        IMAGE_addr <= 5189;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S5206;
      end
      test_b1_S5206: begin
        IMAGE_addr <= 5190;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5203;
        test_state <= test_b1_S5207;
      end
      test_b1_S5207: begin
        IMAGE_addr <= 5191;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 102;
        test_state <= test_b1_S5208;
      end
      test_b1_S5208: begin
        IMAGE_addr <= 5192;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S5209;
      end
      test_b1_S5209: begin
        IMAGE_addr <= 5193;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 110;
        test_state <= test_b1_S5210;
      end
      test_b1_S5210: begin
        IMAGE_addr <= 5194;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 100;
        test_state <= test_b1_S5211;
      end
      test_b1_S5211: begin
        IMAGE_addr <= 5195;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 73;
        test_state <= test_b1_S5212;
      end
      test_b1_S5212: begin
        IMAGE_addr <= 5196;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 110;
        test_state <= test_b1_S5213;
      end
      test_b1_S5213: begin
        IMAGE_addr <= 5197;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 67;
        test_state <= test_b1_S5214;
      end
      test_b1_S5214: begin
        IMAGE_addr <= 5198;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 104;
        test_state <= test_b1_S5215;
      end
      test_b1_S5215: begin
        IMAGE_addr <= 5199;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S5216;
      end
      test_b1_S5216: begin
        IMAGE_addr <= 5200;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S5217;
      end
      test_b1_S5217: begin
        IMAGE_addr <= 5201;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 110;
        test_state <= test_b1_S5218;
      end
      test_b1_S5218: begin
        IMAGE_addr <= 5202;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S5219;
      end
      test_b1_S5219: begin
        IMAGE_addr <= 5203;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S5220;
      end
      test_b1_S5220: begin
        IMAGE_addr <= 5204;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S5221;
      end
      test_b1_S5221: begin
        IMAGE_addr <= 5205;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5116;
        test_state <= test_b1_S5222;
      end
      test_b1_S5222: begin
        IMAGE_addr <= 5206;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1232;
        test_state <= test_b1_S5223;
      end
      test_b1_S5223: begin
        IMAGE_addr <= 5207;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5157;
        test_state <= test_b1_S5224;
      end
      test_b1_S5224: begin
        IMAGE_addr <= 5208;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5225;
      end
      test_b1_S5225: begin
        IMAGE_addr <= 5209;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5226;
      end
      test_b1_S5226: begin
        IMAGE_addr <= 5210;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5188;
        test_state <= test_b1_S5227;
      end
      test_b1_S5227: begin
        IMAGE_addr <= 5211;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S5228;
      end
      test_b1_S5228: begin
        IMAGE_addr <= 5212;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5219;
        test_state <= test_b1_S5229;
      end
      test_b1_S5229: begin
        IMAGE_addr <= 5213;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 119;
        test_state <= test_b1_S5230;
      end
      test_b1_S5230: begin
        IMAGE_addr <= 5214;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S5231;
      end
      test_b1_S5231: begin
        IMAGE_addr <= 5215;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S5232;
      end
      test_b1_S5232: begin
        IMAGE_addr <= 5216;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 104;
        test_state <= test_b1_S5233;
      end
      test_b1_S5233: begin
        IMAGE_addr <= 5217;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 124;
        test_state <= test_b1_S5234;
      end
      test_b1_S5234: begin
        IMAGE_addr <= 5218;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S5235;
      end
      test_b1_S5235: begin
        IMAGE_addr <= 5219;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S5236;
      end
      test_b1_S5236: begin
        IMAGE_addr <= 5220;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S5237;
      end
      test_b1_S5237: begin
        IMAGE_addr <= 5221;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5179;
        test_state <= test_b1_S5238;
      end
      test_b1_S5238: begin
        IMAGE_addr <= 5222;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5239;
      end
      test_b1_S5239: begin
        IMAGE_addr <= 5223;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 32;
        test_state <= test_b1_S5240;
      end
      test_b1_S5240: begin
        IMAGE_addr <= 5224;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 562;
        test_state <= test_b1_S5241;
      end
      test_b1_S5241: begin
        IMAGE_addr <= 5225;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 400;
        test_state <= test_b1_S5242;
      end
      test_b1_S5242: begin
        IMAGE_addr <= 5226;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5243;
      end
      test_b1_S5243: begin
        IMAGE_addr <= 5227;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4905;
        test_state <= test_b1_S5244;
      end
      test_b1_S5244: begin
        IMAGE_addr <= 5228;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 838;
        test_state <= test_b1_S5245;
      end
      test_b1_S5245: begin
        IMAGE_addr <= 5229;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 140;
        test_state <= test_b1_S5246;
      end
      test_b1_S5246: begin
        IMAGE_addr <= 5230;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 25;
        test_state <= test_b1_S5247;
      end
      test_b1_S5247: begin
        IMAGE_addr <= 5231;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S5248;
      end
      test_b1_S5248: begin
        IMAGE_addr <= 5232;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 400;
        test_state <= test_b1_S5249;
      end
      test_b1_S5249: begin
        IMAGE_addr <= 5233;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1232;
        test_state <= test_b1_S5250;
      end
      test_b1_S5250: begin
        IMAGE_addr <= 5234;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S5251;
      end
      test_b1_S5251: begin
        IMAGE_addr <= 5235;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5240;
        test_state <= test_b1_S5252;
      end
      test_b1_S5252: begin
        IMAGE_addr <= 5236;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 583;
        test_state <= test_b1_S5253;
      end
      test_b1_S5253: begin
        IMAGE_addr <= 5237;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S5254;
      end
      test_b1_S5254: begin
        IMAGE_addr <= 5238;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5116;
        test_state <= test_b1_S5255;
      end
      test_b1_S5255: begin
        IMAGE_addr <= 5239;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5256;
      end
      test_b1_S5256: begin
        IMAGE_addr <= 5240;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5257;
      end
      test_b1_S5257: begin
        IMAGE_addr <= 5241;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 52;
        test_state <= test_b1_S5258;
      end
      test_b1_S5258: begin
        IMAGE_addr <= 5242;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 732;
        test_state <= test_b1_S5259;
      end
      test_b1_S5259: begin
        IMAGE_addr <= 5243;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8;
        test_state <= test_b1_S5260;
      end
      test_b1_S5260: begin
        IMAGE_addr <= 5244;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5222;
        test_state <= test_b1_S5261;
      end
      test_b1_S5261: begin
        IMAGE_addr <= 5245;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5262;
      end
      test_b1_S5262: begin
        IMAGE_addr <= 5246;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5263;
      end
      test_b1_S5263: begin
        IMAGE_addr <= 5247;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5210;
        test_state <= test_b1_S5264;
      end
      test_b1_S5264: begin
        IMAGE_addr <= 5248;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S5265;
      end
      test_b1_S5265: begin
        IMAGE_addr <= 5249;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5258;
        test_state <= test_b1_S5266;
      end
      test_b1_S5266: begin
        IMAGE_addr <= 5250;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S5267;
      end
      test_b1_S5267: begin
        IMAGE_addr <= 5251;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S5268;
      end
      test_b1_S5268: begin
        IMAGE_addr <= 5252;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 110;
        test_state <= test_b1_S5269;
      end
      test_b1_S5269: begin
        IMAGE_addr <= 5253;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S5270;
      end
      test_b1_S5270: begin
        IMAGE_addr <= 5254;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 109;
        test_state <= test_b1_S5271;
      end
      test_b1_S5271: begin
        IMAGE_addr <= 5255;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S5272;
      end
      test_b1_S5272: begin
        IMAGE_addr <= 5256;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 58;
        test_state <= test_b1_S5273;
      end
      test_b1_S5273: begin
        IMAGE_addr <= 5257;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S5274;
      end
      test_b1_S5274: begin
        IMAGE_addr <= 5258;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S5275;
      end
      test_b1_S5275: begin
        IMAGE_addr <= 5259;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S5276;
      end
      test_b1_S5276: begin
        IMAGE_addr <= 5260;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 621;
        test_state <= test_b1_S5277;
      end
      test_b1_S5277: begin
        IMAGE_addr <= 5261;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S5278;
      end
      test_b1_S5278: begin
        IMAGE_addr <= 5262;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3056;
        test_state <= test_b1_S5279;
      end
      test_b1_S5279: begin
        IMAGE_addr <= 5263;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S5280;
      end
      test_b1_S5280: begin
        IMAGE_addr <= 5264;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3083;
        test_state <= test_b1_S5281;
      end
      test_b1_S5281: begin
        IMAGE_addr <= 5265;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S5282;
      end
      test_b1_S5282: begin
        IMAGE_addr <= 5266;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5275;
        test_state <= test_b1_S5283;
      end
      test_b1_S5283: begin
        IMAGE_addr <= 5267;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 583;
        test_state <= test_b1_S5284;
      end
      test_b1_S5284: begin
        IMAGE_addr <= 5268;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S5285;
      end
      test_b1_S5285: begin
        IMAGE_addr <= 5269;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5286;
      end
      test_b1_S5286: begin
        IMAGE_addr <= 5270;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S5287;
      end
      test_b1_S5287: begin
        IMAGE_addr <= 5271;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S5288;
      end
      test_b1_S5288: begin
        IMAGE_addr <= 5272;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 583;
        test_state <= test_b1_S5289;
      end
      test_b1_S5289: begin
        IMAGE_addr <= 5273;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S5290;
      end
      test_b1_S5290: begin
        IMAGE_addr <= 5274;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5291;
      end
      test_b1_S5291: begin
        IMAGE_addr <= 5275;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S5292;
      end
      test_b1_S5292: begin
        IMAGE_addr <= 5276;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5285;
        test_state <= test_b1_S5293;
      end
      test_b1_S5293: begin
        IMAGE_addr <= 5277;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 578;
        test_state <= test_b1_S5294;
      end
      test_b1_S5294: begin
        IMAGE_addr <= 5278;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S5295;
      end
      test_b1_S5295: begin
        IMAGE_addr <= 5279;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5296;
      end
      test_b1_S5296: begin
        IMAGE_addr <= 5280;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S5297;
      end
      test_b1_S5297: begin
        IMAGE_addr <= 5281;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S5298;
      end
      test_b1_S5298: begin
        IMAGE_addr <= 5282;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 578;
        test_state <= test_b1_S5299;
      end
      test_b1_S5299: begin
        IMAGE_addr <= 5283;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S5300;
      end
      test_b1_S5300: begin
        IMAGE_addr <= 5284;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5301;
      end
      test_b1_S5301: begin
        IMAGE_addr <= 5285;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3539;
        test_state <= test_b1_S5302;
      end
      test_b1_S5302: begin
        IMAGE_addr <= 5286;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5303;
      end
      test_b1_S5303: begin
        IMAGE_addr <= 5287;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5304;
      end
      test_b1_S5304: begin
        IMAGE_addr <= 5288;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S5305;
      end
      test_b1_S5305: begin
        IMAGE_addr <= 5289;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S5306;
      end
      test_b1_S5306: begin
        IMAGE_addr <= 5290;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2314;
        test_state <= test_b1_S5307;
      end
      test_b1_S5307: begin
        IMAGE_addr <= 5291;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8479;
        test_state <= test_b1_S5308;
      end
      test_b1_S5308: begin
        IMAGE_addr <= 5292;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5421;
        test_state <= test_b1_S5309;
      end
      test_b1_S5309: begin
        IMAGE_addr <= 5293;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5247;
        test_state <= test_b1_S5310;
      end
      test_b1_S5310: begin
        IMAGE_addr <= 5294;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 310;
        test_state <= test_b1_S5311;
      end
      test_b1_S5311: begin
        IMAGE_addr <= 5295;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5288;
        test_state <= test_b1_S5312;
      end
      test_b1_S5312: begin
        IMAGE_addr <= 5296;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 102;
        test_state <= test_b1_S5313;
      end
      test_b1_S5313: begin
        IMAGE_addr <= 5297;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 108;
        test_state <= test_b1_S5314;
      end
      test_b1_S5314: begin
        IMAGE_addr <= 5298;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S5315;
      end
      test_b1_S5315: begin
        IMAGE_addr <= 5299;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 103;
        test_state <= test_b1_S5316;
      end
      test_b1_S5316: begin
        IMAGE_addr <= 5300;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S5317;
      end
      test_b1_S5317: begin
        IMAGE_addr <= 5301;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5293;
        test_state <= test_b1_S5318;
      end
      test_b1_S5318: begin
        IMAGE_addr <= 5302;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 310;
        test_state <= test_b1_S5319;
      end
      test_b1_S5319: begin
        IMAGE_addr <= 5303;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5289;
        test_state <= test_b1_S5320;
      end
      test_b1_S5320: begin
        IMAGE_addr <= 5304;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 100;
        test_state <= test_b1_S5321;
      end
      test_b1_S5321: begin
        IMAGE_addr <= 5305;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S5322;
      end
      test_b1_S5322: begin
        IMAGE_addr <= 5306;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S5323;
      end
      test_b1_S5323: begin
        IMAGE_addr <= 5307;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5301;
        test_state <= test_b1_S5324;
      end
      test_b1_S5324: begin
        IMAGE_addr <= 5308;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 310;
        test_state <= test_b1_S5325;
      end
      test_b1_S5325: begin
        IMAGE_addr <= 5309;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5290;
        test_state <= test_b1_S5326;
      end
      test_b1_S5326: begin
        IMAGE_addr <= 5310;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 110;
        test_state <= test_b1_S5327;
      end
      test_b1_S5327: begin
        IMAGE_addr <= 5311;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S5328;
      end
      test_b1_S5328: begin
        IMAGE_addr <= 5312;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 109;
        test_state <= test_b1_S5329;
      end
      test_b1_S5329: begin
        IMAGE_addr <= 5313;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S5330;
      end
      test_b1_S5330: begin
        IMAGE_addr <= 5314;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S5331;
      end
      test_b1_S5331: begin
        IMAGE_addr <= 5315;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5307;
        test_state <= test_b1_S5332;
      end
      test_b1_S5332: begin
        IMAGE_addr <= 5316;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 310;
        test_state <= test_b1_S5333;
      end
      test_b1_S5333: begin
        IMAGE_addr <= 5317;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5291;
        test_state <= test_b1_S5334;
      end
      test_b1_S5334: begin
        IMAGE_addr <= 5318;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S5335;
      end
      test_b1_S5335: begin
        IMAGE_addr <= 5319;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S5336;
      end
      test_b1_S5336: begin
        IMAGE_addr <= 5320;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 102;
        test_state <= test_b1_S5337;
      end
      test_b1_S5337: begin
        IMAGE_addr <= 5321;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S5338;
      end
      test_b1_S5338: begin
        IMAGE_addr <= 5322;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S5339;
      end
      test_b1_S5339: begin
        IMAGE_addr <= 5323;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 121;
        test_state <= test_b1_S5340;
      end
      test_b1_S5340: begin
        IMAGE_addr <= 5324;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S5341;
      end
      test_b1_S5341: begin
        IMAGE_addr <= 5325;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5315;
        test_state <= test_b1_S5342;
      end
      test_b1_S5342: begin
        IMAGE_addr <= 5326;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 310;
        test_state <= test_b1_S5343;
      end
      test_b1_S5343: begin
        IMAGE_addr <= 5327;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5292;
        test_state <= test_b1_S5344;
      end
      test_b1_S5344: begin
        IMAGE_addr <= 5328;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 120;
        test_state <= test_b1_S5345;
      end
      test_b1_S5345: begin
        IMAGE_addr <= 5329;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S5346;
      end
      test_b1_S5346: begin
        IMAGE_addr <= 5330;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S5347;
      end
      test_b1_S5347: begin
        IMAGE_addr <= 5331;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5325;
        test_state <= test_b1_S5348;
      end
      test_b1_S5348: begin
        IMAGE_addr <= 5332;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S5349;
      end
      test_b1_S5349: begin
        IMAGE_addr <= 5333;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5341;
        test_state <= test_b1_S5350;
      end
      test_b1_S5350: begin
        IMAGE_addr <= 5334;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S5351;
      end
      test_b1_S5351: begin
        IMAGE_addr <= 5335;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S5352;
      end
      test_b1_S5352: begin
        IMAGE_addr <= 5336;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S5353;
      end
      test_b1_S5353: begin
        IMAGE_addr <= 5337;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S5354;
      end
      test_b1_S5354: begin
        IMAGE_addr <= 5338;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 99;
        test_state <= test_b1_S5355;
      end
      test_b1_S5355: begin
        IMAGE_addr <= 5339;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 104;
        test_state <= test_b1_S5356;
      end
      test_b1_S5356: begin
        IMAGE_addr <= 5340;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S5357;
      end
      test_b1_S5357: begin
        IMAGE_addr <= 5341;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5358;
      end
      test_b1_S5358: begin
        IMAGE_addr <= 5342;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4813;
        test_state <= test_b1_S5359;
      end
      test_b1_S5359: begin
        IMAGE_addr <= 5343;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S5360;
      end
      test_b1_S5360: begin
        IMAGE_addr <= 5344;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 25;
        test_state <= test_b1_S5361;
      end
      test_b1_S5361: begin
        IMAGE_addr <= 5345;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S5362;
      end
      test_b1_S5362: begin
        IMAGE_addr <= 5346;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5363;
      end
      test_b1_S5363: begin
        IMAGE_addr <= 5347;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4813;
        test_state <= test_b1_S5364;
      end
      test_b1_S5364: begin
        IMAGE_addr <= 5348;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 16;
        test_state <= test_b1_S5365;
      end
      test_b1_S5365: begin
        IMAGE_addr <= 5349;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5011;
        test_state <= test_b1_S5366;
      end
      test_b1_S5366: begin
        IMAGE_addr <= 5350;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5367;
      end
      test_b1_S5367: begin
        IMAGE_addr <= 5351;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5292;
        test_state <= test_b1_S5368;
      end
      test_b1_S5368: begin
        IMAGE_addr <= 5352;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S5369;
      end
      test_b1_S5369: begin
        IMAGE_addr <= 5353;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 183;
        test_state <= test_b1_S5370;
      end
      test_b1_S5370: begin
        IMAGE_addr <= 5354;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 27;
        test_state <= test_b1_S5371;
      end
      test_b1_S5371: begin
        IMAGE_addr <= 5355;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8;
        test_state <= test_b1_S5372;
      end
      test_b1_S5372: begin
        IMAGE_addr <= 5356;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5344;
        test_state <= test_b1_S5373;
      end
      test_b1_S5373: begin
        IMAGE_addr <= 5357;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5374;
      end
      test_b1_S5374: begin
        IMAGE_addr <= 5358;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5375;
      end
      test_b1_S5375: begin
        IMAGE_addr <= 5359;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5331;
        test_state <= test_b1_S5376;
      end
      test_b1_S5376: begin
        IMAGE_addr <= 5360;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S5377;
      end
      test_b1_S5377: begin
        IMAGE_addr <= 5361;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5370;
        test_state <= test_b1_S5378;
      end
      test_b1_S5378: begin
        IMAGE_addr <= 5362;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 40;
        test_state <= test_b1_S5379;
      end
      test_b1_S5379: begin
        IMAGE_addr <= 5363;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 99;
        test_state <= test_b1_S5380;
      end
      test_b1_S5380: begin
        IMAGE_addr <= 5364;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 104;
        test_state <= test_b1_S5381;
      end
      test_b1_S5381: begin
        IMAGE_addr <= 5365;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S5382;
      end
      test_b1_S5382: begin
        IMAGE_addr <= 5366;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S5383;
      end
      test_b1_S5383: begin
        IMAGE_addr <= 5367;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 110;
        test_state <= test_b1_S5384;
      end
      test_b1_S5384: begin
        IMAGE_addr <= 5368;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S5385;
      end
      test_b1_S5385: begin
        IMAGE_addr <= 5369;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S5386;
      end
      test_b1_S5386: begin
        IMAGE_addr <= 5370;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5387;
      end
      test_b1_S5387: begin
        IMAGE_addr <= 5371;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5290;
        test_state <= test_b1_S5388;
      end
      test_b1_S5388: begin
        IMAGE_addr <= 5372;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S5389;
      end
      test_b1_S5389: begin
        IMAGE_addr <= 5373;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5390;
      end
      test_b1_S5390: begin
        IMAGE_addr <= 5374;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S5391;
      end
      test_b1_S5391: begin
        IMAGE_addr <= 5375;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S5392;
      end
      test_b1_S5392: begin
        IMAGE_addr <= 5376;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5381;
        test_state <= test_b1_S5393;
      end
      test_b1_S5393: begin
        IMAGE_addr <= 5377;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5394;
      end
      test_b1_S5394: begin
        IMAGE_addr <= 5378;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5289;
        test_state <= test_b1_S5395;
      end
      test_b1_S5395: begin
        IMAGE_addr <= 5379;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S5396;
      end
      test_b1_S5396: begin
        IMAGE_addr <= 5380;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5397;
      end
      test_b1_S5397: begin
        IMAGE_addr <= 5381;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S5398;
      end
      test_b1_S5398: begin
        IMAGE_addr <= 5382;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5387;
        test_state <= test_b1_S5399;
      end
      test_b1_S5399: begin
        IMAGE_addr <= 5383;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5400;
      end
      test_b1_S5400: begin
        IMAGE_addr <= 5384;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5288;
        test_state <= test_b1_S5401;
      end
      test_b1_S5401: begin
        IMAGE_addr <= 5385;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S5402;
      end
      test_b1_S5402: begin
        IMAGE_addr <= 5386;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5403;
      end
      test_b1_S5403: begin
        IMAGE_addr <= 5387;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3539;
        test_state <= test_b1_S5404;
      end
      test_b1_S5404: begin
        IMAGE_addr <= 5388;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5405;
      end
      test_b1_S5405: begin
        IMAGE_addr <= 5389;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S5406;
      end
      test_b1_S5406: begin
        IMAGE_addr <= 5390;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S5407;
      end
      test_b1_S5407: begin
        IMAGE_addr <= 5391;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5408;
      end
      test_b1_S5408: begin
        IMAGE_addr <= 5392;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5291;
        test_state <= test_b1_S5409;
      end
      test_b1_S5409: begin
        IMAGE_addr <= 5393;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S5410;
      end
      test_b1_S5410: begin
        IMAGE_addr <= 5394;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5411;
      end
      test_b1_S5411: begin
        IMAGE_addr <= 5395;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5412;
      end
      test_b1_S5412: begin
        IMAGE_addr <= 5396;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5359;
        test_state <= test_b1_S5413;
      end
      test_b1_S5413: begin
        IMAGE_addr <= 5397;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S5414;
      end
      test_b1_S5414: begin
        IMAGE_addr <= 5398;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5405;
        test_state <= test_b1_S5415;
      end
      test_b1_S5415: begin
        IMAGE_addr <= 5399;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 98;
        test_state <= test_b1_S5416;
      end
      test_b1_S5416: begin
        IMAGE_addr <= 5400;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S5417;
      end
      test_b1_S5417: begin
        IMAGE_addr <= 5401;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 99;
        test_state <= test_b1_S5418;
      end
      test_b1_S5418: begin
        IMAGE_addr <= 5402;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 107;
        test_state <= test_b1_S5419;
      end
      test_b1_S5419: begin
        IMAGE_addr <= 5403;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 41;
        test_state <= test_b1_S5420;
      end
      test_b1_S5420: begin
        IMAGE_addr <= 5404;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S5421;
      end
      test_b1_S5421: begin
        IMAGE_addr <= 5405;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5422;
      end
      test_b1_S5422: begin
        IMAGE_addr <= 5406;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5291;
        test_state <= test_b1_S5423;
      end
      test_b1_S5423: begin
        IMAGE_addr <= 5407;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S5424;
      end
      test_b1_S5424: begin
        IMAGE_addr <= 5408;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5425;
      end
      test_b1_S5425: begin
        IMAGE_addr <= 5409;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S5426;
      end
      test_b1_S5426: begin
        IMAGE_addr <= 5410;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S5427;
      end
      test_b1_S5427: begin
        IMAGE_addr <= 5411;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5428;
      end
      test_b1_S5428: begin
        IMAGE_addr <= 5412;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5429;
      end
      test_b1_S5429: begin
        IMAGE_addr <= 5413;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5396;
        test_state <= test_b1_S5430;
      end
      test_b1_S5430: begin
        IMAGE_addr <= 5414;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S5431;
      end
      test_b1_S5431: begin
        IMAGE_addr <= 5415;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5421;
        test_state <= test_b1_S5432;
      end
      test_b1_S5432: begin
        IMAGE_addr <= 5416;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S5433;
      end
      test_b1_S5433: begin
        IMAGE_addr <= 5417;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S5434;
      end
      test_b1_S5434: begin
        IMAGE_addr <= 5418;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S5435;
      end
      test_b1_S5435: begin
        IMAGE_addr <= 5419;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 107;
        test_state <= test_b1_S5436;
      end
      test_b1_S5436: begin
        IMAGE_addr <= 5420;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S5437;
      end
      test_b1_S5437: begin
        IMAGE_addr <= 5421;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5438;
      end
      test_b1_S5438: begin
        IMAGE_addr <= 5422;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5290;
        test_state <= test_b1_S5439;
      end
      test_b1_S5439: begin
        IMAGE_addr <= 5423;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S5440;
      end
      test_b1_S5440: begin
        IMAGE_addr <= 5424;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1234;
        test_state <= test_b1_S5441;
      end
      test_b1_S5441: begin
        IMAGE_addr <= 5425;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S5442;
      end
      test_b1_S5442: begin
        IMAGE_addr <= 5426;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5437;
        test_state <= test_b1_S5443;
      end
      test_b1_S5443: begin
        IMAGE_addr <= 5427;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5444;
      end
      test_b1_S5444: begin
        IMAGE_addr <= 5428;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5289;
        test_state <= test_b1_S5445;
      end
      test_b1_S5445: begin
        IMAGE_addr <= 5429;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S5446;
      end
      test_b1_S5446: begin
        IMAGE_addr <= 5430;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5447;
      end
      test_b1_S5447: begin
        IMAGE_addr <= 5431;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5288;
        test_state <= test_b1_S5448;
      end
      test_b1_S5448: begin
        IMAGE_addr <= 5432;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 147;
        test_state <= test_b1_S5449;
      end
      test_b1_S5449: begin
        IMAGE_addr <= 5433;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S5450;
      end
      test_b1_S5450: begin
        IMAGE_addr <= 5434;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5451;
      end
      test_b1_S5451: begin
        IMAGE_addr <= 5435;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5452;
      end
      test_b1_S5452: begin
        IMAGE_addr <= 5436;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5453;
      end
      test_b1_S5453: begin
        IMAGE_addr <= 5437;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5454;
      end
      test_b1_S5454: begin
        IMAGE_addr <= 5438;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 52;
        test_state <= test_b1_S5455;
      end
      test_b1_S5455: begin
        IMAGE_addr <= 5439;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 732;
        test_state <= test_b1_S5456;
      end
      test_b1_S5456: begin
        IMAGE_addr <= 5440;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5457;
      end
      test_b1_S5457: begin
        IMAGE_addr <= 5441;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5458;
      end
      test_b1_S5458: begin
        IMAGE_addr <= 5442;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5413;
        test_state <= test_b1_S5459;
      end
      test_b1_S5459: begin
        IMAGE_addr <= 5443;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S5460;
      end
      test_b1_S5460: begin
        IMAGE_addr <= 5444;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5452;
        test_state <= test_b1_S5461;
      end
      test_b1_S5461: begin
        IMAGE_addr <= 5445;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 108;
        test_state <= test_b1_S5462;
      end
      test_b1_S5462: begin
        IMAGE_addr <= 5446;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 111;
        test_state <= test_b1_S5463;
      end
      test_b1_S5463: begin
        IMAGE_addr <= 5447;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 111;
        test_state <= test_b1_S5464;
      end
      test_b1_S5464: begin
        IMAGE_addr <= 5448;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 107;
        test_state <= test_b1_S5465;
      end
      test_b1_S5465: begin
        IMAGE_addr <= 5449;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 117;
        test_state <= test_b1_S5466;
      end
      test_b1_S5466: begin
        IMAGE_addr <= 5450;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 112;
        test_state <= test_b1_S5467;
      end
      test_b1_S5467: begin
        IMAGE_addr <= 5451;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S5468;
      end
      test_b1_S5468: begin
        IMAGE_addr <= 5452;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5469;
      end
      test_b1_S5469: begin
        IMAGE_addr <= 5453;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5421;
        test_state <= test_b1_S5470;
      end
      test_b1_S5470: begin
        IMAGE_addr <= 5454;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5471;
      end
      test_b1_S5471: begin
        IMAGE_addr <= 5455;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5292;
        test_state <= test_b1_S5472;
      end
      test_b1_S5472: begin
        IMAGE_addr <= 5456;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S5473;
      end
      test_b1_S5473: begin
        IMAGE_addr <= 5457;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5370;
        test_state <= test_b1_S5474;
      end
      test_b1_S5474: begin
        IMAGE_addr <= 5458;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5341;
        test_state <= test_b1_S5475;
      end
      test_b1_S5475: begin
        IMAGE_addr <= 5459;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5405;
        test_state <= test_b1_S5476;
      end
      test_b1_S5476: begin
        IMAGE_addr <= 5460;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5477;
      end
      test_b1_S5477: begin
        IMAGE_addr <= 5461;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5288;
        test_state <= test_b1_S5478;
      end
      test_b1_S5478: begin
        IMAGE_addr <= 5462;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S5479;
      end
      test_b1_S5479: begin
        IMAGE_addr <= 5463;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S5480;
      end
      test_b1_S5480: begin
        IMAGE_addr <= 5464;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5472;
        test_state <= test_b1_S5481;
      end
      test_b1_S5481: begin
        IMAGE_addr <= 5465;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5482;
      end
      test_b1_S5482: begin
        IMAGE_addr <= 5466;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5289;
        test_state <= test_b1_S5483;
      end
      test_b1_S5483: begin
        IMAGE_addr <= 5467;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S5484;
      end
      test_b1_S5484: begin
        IMAGE_addr <= 5468;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5485;
      end
      test_b1_S5485: begin
        IMAGE_addr <= 5469;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5288;
        test_state <= test_b1_S5486;
      end
      test_b1_S5486: begin
        IMAGE_addr <= 5470;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S5487;
      end
      test_b1_S5487: begin
        IMAGE_addr <= 5471;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5488;
      end
      test_b1_S5488: begin
        IMAGE_addr <= 5472;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S5489;
      end
      test_b1_S5489: begin
        IMAGE_addr <= 5473;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5479;
        test_state <= test_b1_S5490;
      end
      test_b1_S5490: begin
        IMAGE_addr <= 5474;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5491;
      end
      test_b1_S5491: begin
        IMAGE_addr <= 5475;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5290;
        test_state <= test_b1_S5492;
      end
      test_b1_S5492: begin
        IMAGE_addr <= 5476;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S5493;
      end
      test_b1_S5493: begin
        IMAGE_addr <= 5477;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1234;
        test_state <= test_b1_S5494;
      end
      test_b1_S5494: begin
        IMAGE_addr <= 5478;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5495;
      end
      test_b1_S5495: begin
        IMAGE_addr <= 5479;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 732;
        test_state <= test_b1_S5496;
      end
      test_b1_S5496: begin
        IMAGE_addr <= 5480;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5497;
      end
      test_b1_S5497: begin
        IMAGE_addr <= 5481;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5498;
      end
      test_b1_S5498: begin
        IMAGE_addr <= 5482;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5442;
        test_state <= test_b1_S5499;
      end
      test_b1_S5499: begin
        IMAGE_addr <= 5483;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S5500;
      end
      test_b1_S5500: begin
        IMAGE_addr <= 5484;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5490;
        test_state <= test_b1_S5501;
      end
      test_b1_S5501: begin
        IMAGE_addr <= 5485;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S5502;
      end
      test_b1_S5502: begin
        IMAGE_addr <= 5486;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S5503;
      end
      test_b1_S5503: begin
        IMAGE_addr <= 5487;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S5504;
      end
      test_b1_S5504: begin
        IMAGE_addr <= 5488;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 107;
        test_state <= test_b1_S5505;
      end
      test_b1_S5505: begin
        IMAGE_addr <= 5489;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S5506;
      end
      test_b1_S5506: begin
        IMAGE_addr <= 5490;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5507;
      end
      test_b1_S5507: begin
        IMAGE_addr <= 5491;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5290;
        test_state <= test_b1_S5508;
      end
      test_b1_S5508: begin
        IMAGE_addr <= 5492;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S5509;
      end
      test_b1_S5509: begin
        IMAGE_addr <= 5493;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3058;
        test_state <= test_b1_S5510;
      end
      test_b1_S5510: begin
        IMAGE_addr <= 5494;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S5511;
      end
      test_b1_S5511: begin
        IMAGE_addr <= 5495;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S5512;
      end
      test_b1_S5512: begin
        IMAGE_addr <= 5496;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5507;
        test_state <= test_b1_S5513;
      end
      test_b1_S5513: begin
        IMAGE_addr <= 5497;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5514;
      end
      test_b1_S5514: begin
        IMAGE_addr <= 5498;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5289;
        test_state <= test_b1_S5515;
      end
      test_b1_S5515: begin
        IMAGE_addr <= 5499;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S5516;
      end
      test_b1_S5516: begin
        IMAGE_addr <= 5500;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5517;
      end
      test_b1_S5517: begin
        IMAGE_addr <= 5501;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5288;
        test_state <= test_b1_S5518;
      end
      test_b1_S5518: begin
        IMAGE_addr <= 5502;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 147;
        test_state <= test_b1_S5519;
      end
      test_b1_S5519: begin
        IMAGE_addr <= 5503;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S5520;
      end
      test_b1_S5520: begin
        IMAGE_addr <= 5504;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5521;
      end
      test_b1_S5521: begin
        IMAGE_addr <= 5505;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5522;
      end
      test_b1_S5522: begin
        IMAGE_addr <= 5506;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5523;
      end
      test_b1_S5523: begin
        IMAGE_addr <= 5507;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5524;
      end
      test_b1_S5524: begin
        IMAGE_addr <= 5508;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 52;
        test_state <= test_b1_S5525;
      end
      test_b1_S5525: begin
        IMAGE_addr <= 5509;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 732;
        test_state <= test_b1_S5526;
      end
      test_b1_S5526: begin
        IMAGE_addr <= 5510;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5527;
      end
      test_b1_S5527: begin
        IMAGE_addr <= 5511;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5528;
      end
      test_b1_S5528: begin
        IMAGE_addr <= 5512;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5482;
        test_state <= test_b1_S5529;
      end
      test_b1_S5529: begin
        IMAGE_addr <= 5513;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S5530;
      end
      test_b1_S5530: begin
        IMAGE_addr <= 5514;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5522;
        test_state <= test_b1_S5531;
      end
      test_b1_S5531: begin
        IMAGE_addr <= 5515;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 108;
        test_state <= test_b1_S5532;
      end
      test_b1_S5532: begin
        IMAGE_addr <= 5516;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 111;
        test_state <= test_b1_S5533;
      end
      test_b1_S5533: begin
        IMAGE_addr <= 5517;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 111;
        test_state <= test_b1_S5534;
      end
      test_b1_S5534: begin
        IMAGE_addr <= 5518;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 107;
        test_state <= test_b1_S5535;
      end
      test_b1_S5535: begin
        IMAGE_addr <= 5519;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 117;
        test_state <= test_b1_S5536;
      end
      test_b1_S5536: begin
        IMAGE_addr <= 5520;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 112;
        test_state <= test_b1_S5537;
      end
      test_b1_S5537: begin
        IMAGE_addr <= 5521;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S5538;
      end
      test_b1_S5538: begin
        IMAGE_addr <= 5522;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5539;
      end
      test_b1_S5539: begin
        IMAGE_addr <= 5523;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5490;
        test_state <= test_b1_S5540;
      end
      test_b1_S5540: begin
        IMAGE_addr <= 5524;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5541;
      end
      test_b1_S5541: begin
        IMAGE_addr <= 5525;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5292;
        test_state <= test_b1_S5542;
      end
      test_b1_S5542: begin
        IMAGE_addr <= 5526;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S5543;
      end
      test_b1_S5543: begin
        IMAGE_addr <= 5527;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5370;
        test_state <= test_b1_S5544;
      end
      test_b1_S5544: begin
        IMAGE_addr <= 5528;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5341;
        test_state <= test_b1_S5545;
      end
      test_b1_S5545: begin
        IMAGE_addr <= 5529;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5405;
        test_state <= test_b1_S5546;
      end
      test_b1_S5546: begin
        IMAGE_addr <= 5530;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5547;
      end
      test_b1_S5547: begin
        IMAGE_addr <= 5531;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5288;
        test_state <= test_b1_S5548;
      end
      test_b1_S5548: begin
        IMAGE_addr <= 5532;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S5549;
      end
      test_b1_S5549: begin
        IMAGE_addr <= 5533;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S5550;
      end
      test_b1_S5550: begin
        IMAGE_addr <= 5534;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5539;
        test_state <= test_b1_S5551;
      end
      test_b1_S5551: begin
        IMAGE_addr <= 5535;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5552;
      end
      test_b1_S5552: begin
        IMAGE_addr <= 5536;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5289;
        test_state <= test_b1_S5553;
      end
      test_b1_S5553: begin
        IMAGE_addr <= 5537;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S5554;
      end
      test_b1_S5554: begin
        IMAGE_addr <= 5538;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5555;
      end
      test_b1_S5555: begin
        IMAGE_addr <= 5539;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S5556;
      end
      test_b1_S5556: begin
        IMAGE_addr <= 5540;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5546;
        test_state <= test_b1_S5557;
      end
      test_b1_S5557: begin
        IMAGE_addr <= 5541;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5558;
      end
      test_b1_S5558: begin
        IMAGE_addr <= 5542;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5290;
        test_state <= test_b1_S5559;
      end
      test_b1_S5559: begin
        IMAGE_addr <= 5543;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S5560;
      end
      test_b1_S5560: begin
        IMAGE_addr <= 5544;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3058;
        test_state <= test_b1_S5561;
      end
      test_b1_S5561: begin
        IMAGE_addr <= 5545;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5562;
      end
      test_b1_S5562: begin
        IMAGE_addr <= 5546;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 732;
        test_state <= test_b1_S5563;
      end
      test_b1_S5563: begin
        IMAGE_addr <= 5547;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5564;
      end
      test_b1_S5564: begin
        IMAGE_addr <= 5548;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5565;
      end
      test_b1_S5565: begin
        IMAGE_addr <= 5549;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3202;
        test_state <= test_b1_S5566;
      end
      test_b1_S5566: begin
        IMAGE_addr <= 5550;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 306;
        test_state <= test_b1_S5567;
      end
      test_b1_S5567: begin
        IMAGE_addr <= 5551;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2315;
        test_state <= test_b1_S5568;
      end
      test_b1_S5568: begin
        IMAGE_addr <= 5552;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S5569;
      end
      test_b1_S5569: begin
        IMAGE_addr <= 5553;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5247;
        test_state <= test_b1_S5570;
      end
      test_b1_S5570: begin
        IMAGE_addr <= 5554;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 310;
        test_state <= test_b1_S5571;
      end
      test_b1_S5571: begin
        IMAGE_addr <= 5555;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5549;
        test_state <= test_b1_S5572;
      end
      test_b1_S5572: begin
        IMAGE_addr <= 5556;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 120;
        test_state <= test_b1_S5573;
      end
      test_b1_S5573: begin
        IMAGE_addr <= 5557;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S5574;
      end
      test_b1_S5574: begin
        IMAGE_addr <= 5558;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S5575;
      end
      test_b1_S5575: begin
        IMAGE_addr <= 5559;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5553;
        test_state <= test_b1_S5576;
      end
      test_b1_S5576: begin
        IMAGE_addr <= 5560;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 310;
        test_state <= test_b1_S5577;
      end
      test_b1_S5577: begin
        IMAGE_addr <= 5561;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5550;
        test_state <= test_b1_S5578;
      end
      test_b1_S5578: begin
        IMAGE_addr <= 5562;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 99;
        test_state <= test_b1_S5579;
      end
      test_b1_S5579: begin
        IMAGE_addr <= 5563;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 108;
        test_state <= test_b1_S5580;
      end
      test_b1_S5580: begin
        IMAGE_addr <= 5564;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S5581;
      end
      test_b1_S5581: begin
        IMAGE_addr <= 5565;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S5582;
      end
      test_b1_S5582: begin
        IMAGE_addr <= 5566;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S5583;
      end
      test_b1_S5583: begin
        IMAGE_addr <= 5567;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S5584;
      end
      test_b1_S5584: begin
        IMAGE_addr <= 5568;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5559;
        test_state <= test_b1_S5585;
      end
      test_b1_S5585: begin
        IMAGE_addr <= 5569;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 310;
        test_state <= test_b1_S5586;
      end
      test_b1_S5586: begin
        IMAGE_addr <= 5570;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5551;
        test_state <= test_b1_S5587;
      end
      test_b1_S5587: begin
        IMAGE_addr <= 5571;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 110;
        test_state <= test_b1_S5588;
      end
      test_b1_S5588: begin
        IMAGE_addr <= 5572;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S5589;
      end
      test_b1_S5589: begin
        IMAGE_addr <= 5573;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 109;
        test_state <= test_b1_S5590;
      end
      test_b1_S5590: begin
        IMAGE_addr <= 5574;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S5591;
      end
      test_b1_S5591: begin
        IMAGE_addr <= 5575;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S5592;
      end
      test_b1_S5592: begin
        IMAGE_addr <= 5576;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5568;
        test_state <= test_b1_S5593;
      end
      test_b1_S5593: begin
        IMAGE_addr <= 5577;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 310;
        test_state <= test_b1_S5594;
      end
      test_b1_S5594: begin
        IMAGE_addr <= 5578;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5552;
        test_state <= test_b1_S5595;
      end
      test_b1_S5595: begin
        IMAGE_addr <= 5579;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 102;
        test_state <= test_b1_S5596;
      end
      test_b1_S5596: begin
        IMAGE_addr <= 5580;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 108;
        test_state <= test_b1_S5597;
      end
      test_b1_S5597: begin
        IMAGE_addr <= 5581;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S5598;
      end
      test_b1_S5598: begin
        IMAGE_addr <= 5582;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 103;
        test_state <= test_b1_S5599;
      end
      test_b1_S5599: begin
        IMAGE_addr <= 5583;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S5600;
      end
      test_b1_S5600: begin
        IMAGE_addr <= 5584;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5576;
        test_state <= test_b1_S5601;
      end
      test_b1_S5601: begin
        IMAGE_addr <= 5585;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 310;
        test_state <= test_b1_S5602;
      end
      test_b1_S5602: begin
        IMAGE_addr <= 5586;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5591;
        test_state <= test_b1_S5603;
      end
      test_b1_S5603: begin
        IMAGE_addr <= 5587;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 95;
        test_state <= test_b1_S5604;
      end
      test_b1_S5604: begin
        IMAGE_addr <= 5588;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 95;
        test_state <= test_b1_S5605;
      end
      test_b1_S5605: begin
        IMAGE_addr <= 5589;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 95;
        test_state <= test_b1_S5606;
      end
      test_b1_S5606: begin
        IMAGE_addr <= 5590;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S5607;
      end
      test_b1_S5607: begin
        IMAGE_addr <= 5591;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 95;
        test_state <= test_b1_S5608;
      end
      test_b1_S5608: begin
        IMAGE_addr <= 5592;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 95;
        test_state <= test_b1_S5609;
      end
      test_b1_S5609: begin
        IMAGE_addr <= 5593;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 64;
        test_state <= test_b1_S5610;
      end
      test_b1_S5610: begin
        IMAGE_addr <= 5594;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S5611;
      end
      test_b1_S5611: begin
        IMAGE_addr <= 5595;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5584;
        test_state <= test_b1_S5612;
      end
      test_b1_S5612: begin
        IMAGE_addr <= 5596;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S5613;
      end
      test_b1_S5613: begin
        IMAGE_addr <= 5597;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5605;
        test_state <= test_b1_S5614;
      end
      test_b1_S5614: begin
        IMAGE_addr <= 5598;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S5615;
      end
      test_b1_S5615: begin
        IMAGE_addr <= 5599;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 99;
        test_state <= test_b1_S5616;
      end
      test_b1_S5616: begin
        IMAGE_addr <= 5600;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S5617;
      end
      test_b1_S5617: begin
        IMAGE_addr <= 5601;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S5618;
      end
      test_b1_S5618: begin
        IMAGE_addr <= 5602;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 111;
        test_state <= test_b1_S5619;
      end
      test_b1_S5619: begin
        IMAGE_addr <= 5603;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 110;
        test_state <= test_b1_S5620;
      end
      test_b1_S5620: begin
        IMAGE_addr <= 5604;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S5621;
      end
      test_b1_S5621: begin
        IMAGE_addr <= 5605;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5622;
      end
      test_b1_S5622: begin
        IMAGE_addr <= 5606;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5549;
        test_state <= test_b1_S5623;
      end
      test_b1_S5623: begin
        IMAGE_addr <= 5607;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S5624;
      end
      test_b1_S5624: begin
        IMAGE_addr <= 5608;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5625;
      end
      test_b1_S5625: begin
        IMAGE_addr <= 5609;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5550;
        test_state <= test_b1_S5626;
      end
      test_b1_S5626: begin
        IMAGE_addr <= 5610;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S5627;
      end
      test_b1_S5627: begin
        IMAGE_addr <= 5611;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 286;
        test_state <= test_b1_S5628;
      end
      test_b1_S5628: begin
        IMAGE_addr <= 5612;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5629;
      end
      test_b1_S5629: begin
        IMAGE_addr <= 5613;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5630;
      end
      test_b1_S5630: begin
        IMAGE_addr <= 5614;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5595;
        test_state <= test_b1_S5631;
      end
      test_b1_S5631: begin
        IMAGE_addr <= 5615;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S5632;
      end
      test_b1_S5632: begin
        IMAGE_addr <= 5616;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5624;
        test_state <= test_b1_S5633;
      end
      test_b1_S5633: begin
        IMAGE_addr <= 5617;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 40;
        test_state <= test_b1_S5634;
      end
      test_b1_S5634: begin
        IMAGE_addr <= 5618;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S5635;
      end
      test_b1_S5635: begin
        IMAGE_addr <= 5619;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 112;
        test_state <= test_b1_S5636;
      end
      test_b1_S5636: begin
        IMAGE_addr <= 5620;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 108;
        test_state <= test_b1_S5637;
      end
      test_b1_S5637: begin
        IMAGE_addr <= 5621;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S5638;
      end
      test_b1_S5638: begin
        IMAGE_addr <= 5622;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S5639;
      end
      test_b1_S5639: begin
        IMAGE_addr <= 5623;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S5640;
      end
      test_b1_S5640: begin
        IMAGE_addr <= 5624;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 189;
        test_state <= test_b1_S5641;
      end
      test_b1_S5641: begin
        IMAGE_addr <= 5625;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5642;
      end
      test_b1_S5642: begin
        IMAGE_addr <= 5626;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5591;
        test_state <= test_b1_S5643;
      end
      test_b1_S5643: begin
        IMAGE_addr <= 5627;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2606;
        test_state <= test_b1_S5644;
      end
      test_b1_S5644: begin
        IMAGE_addr <= 5628;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 26;
        test_state <= test_b1_S5645;
      end
      test_b1_S5645: begin
        IMAGE_addr <= 5629;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 26;
        test_state <= test_b1_S5646;
      end
      test_b1_S5646: begin
        IMAGE_addr <= 5630;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S5647;
      end
      test_b1_S5647: begin
        IMAGE_addr <= 5631;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S5648;
      end
      test_b1_S5648: begin
        IMAGE_addr <= 5632;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5649;
      end
      test_b1_S5649: begin
        IMAGE_addr <= 5633;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5551;
        test_state <= test_b1_S5650;
      end
      test_b1_S5650: begin
        IMAGE_addr <= 5634;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S5651;
      end
      test_b1_S5651: begin
        IMAGE_addr <= 5635;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5652;
      end
      test_b1_S5652: begin
        IMAGE_addr <= 5636;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5653;
      end
      test_b1_S5653: begin
        IMAGE_addr <= 5637;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5614;
        test_state <= test_b1_S5654;
      end
      test_b1_S5654: begin
        IMAGE_addr <= 5638;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S5655;
      end
      test_b1_S5655: begin
        IMAGE_addr <= 5639;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5648;
        test_state <= test_b1_S5656;
      end
      test_b1_S5656: begin
        IMAGE_addr <= 5640;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 112;
        test_state <= test_b1_S5657;
      end
      test_b1_S5657: begin
        IMAGE_addr <= 5641;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S5658;
      end
      test_b1_S5658: begin
        IMAGE_addr <= 5642;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S5659;
      end
      test_b1_S5659: begin
        IMAGE_addr <= 5643;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 102;
        test_state <= test_b1_S5660;
      end
      test_b1_S5660: begin
        IMAGE_addr <= 5644;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S5661;
      end
      test_b1_S5661: begin
        IMAGE_addr <= 5645;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 120;
        test_state <= test_b1_S5662;
      end
      test_b1_S5662: begin
        IMAGE_addr <= 5646;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 41;
        test_state <= test_b1_S5663;
      end
      test_b1_S5663: begin
        IMAGE_addr <= 5647;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S5664;
      end
      test_b1_S5664: begin
        IMAGE_addr <= 5648;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1232;
        test_state <= test_b1_S5665;
      end
      test_b1_S5665: begin
        IMAGE_addr <= 5649;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S5666;
      end
      test_b1_S5666: begin
        IMAGE_addr <= 5650;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5671;
        test_state <= test_b1_S5667;
      end
      test_b1_S5667: begin
        IMAGE_addr <= 5651;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S5668;
      end
      test_b1_S5668: begin
        IMAGE_addr <= 5652;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5659;
        test_state <= test_b1_S5669;
      end
      test_b1_S5669: begin
        IMAGE_addr <= 5653;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 578;
        test_state <= test_b1_S5670;
      end
      test_b1_S5670: begin
        IMAGE_addr <= 5654;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S5671;
      end
      test_b1_S5671: begin
        IMAGE_addr <= 5655;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5672;
      end
      test_b1_S5672: begin
        IMAGE_addr <= 5656;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5550;
        test_state <= test_b1_S5673;
      end
      test_b1_S5673: begin
        IMAGE_addr <= 5657;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S5674;
      end
      test_b1_S5674: begin
        IMAGE_addr <= 5658;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5675;
      end
      test_b1_S5675: begin
        IMAGE_addr <= 5659;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S5676;
      end
      test_b1_S5676: begin
        IMAGE_addr <= 5660;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5667;
        test_state <= test_b1_S5677;
      end
      test_b1_S5677: begin
        IMAGE_addr <= 5661;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 583;
        test_state <= test_b1_S5678;
      end
      test_b1_S5678: begin
        IMAGE_addr <= 5662;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S5679;
      end
      test_b1_S5679: begin
        IMAGE_addr <= 5663;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5680;
      end
      test_b1_S5680: begin
        IMAGE_addr <= 5664;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5549;
        test_state <= test_b1_S5681;
      end
      test_b1_S5681: begin
        IMAGE_addr <= 5665;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S5682;
      end
      test_b1_S5682: begin
        IMAGE_addr <= 5666;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5683;
      end
      test_b1_S5683: begin
        IMAGE_addr <= 5667;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3539;
        test_state <= test_b1_S5684;
      end
      test_b1_S5684: begin
        IMAGE_addr <= 5668;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5685;
      end
      test_b1_S5685: begin
        IMAGE_addr <= 5669;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4294967295;
        test_state <= test_b1_S5686;
      end
      test_b1_S5686: begin
        IMAGE_addr <= 5670;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5687;
      end
      test_b1_S5687: begin
        IMAGE_addr <= 5671;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S5688;
      end
      test_b1_S5688: begin
        IMAGE_addr <= 5672;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5676;
        test_state <= test_b1_S5689;
      end
      test_b1_S5689: begin
        IMAGE_addr <= 5673;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5690;
      end
      test_b1_S5690: begin
        IMAGE_addr <= 5674;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S5691;
      end
      test_b1_S5691: begin
        IMAGE_addr <= 5675;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5692;
      end
      test_b1_S5692: begin
        IMAGE_addr <= 5676;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 732;
        test_state <= test_b1_S5693;
      end
      test_b1_S5693: begin
        IMAGE_addr <= 5677;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5694;
      end
      test_b1_S5694: begin
        IMAGE_addr <= 5678;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5695;
      end
      test_b1_S5695: begin
        IMAGE_addr <= 5679;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5637;
        test_state <= test_b1_S5696;
      end
      test_b1_S5696: begin
        IMAGE_addr <= 5680;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S5697;
      end
      test_b1_S5697: begin
        IMAGE_addr <= 5681;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5689;
        test_state <= test_b1_S5698;
      end
      test_b1_S5698: begin
        IMAGE_addr <= 5682;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 104;
        test_state <= test_b1_S5699;
      end
      test_b1_S5699: begin
        IMAGE_addr <= 5683;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S5700;
      end
      test_b1_S5700: begin
        IMAGE_addr <= 5684;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 110;
        test_state <= test_b1_S5701;
      end
      test_b1_S5701: begin
        IMAGE_addr <= 5685;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 100;
        test_state <= test_b1_S5702;
      end
      test_b1_S5702: begin
        IMAGE_addr <= 5686;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 108;
        test_state <= test_b1_S5703;
      end
      test_b1_S5703: begin
        IMAGE_addr <= 5687;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S5704;
      end
      test_b1_S5704: begin
        IMAGE_addr <= 5688;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S5705;
      end
      test_b1_S5705: begin
        IMAGE_addr <= 5689;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5706;
      end
      test_b1_S5706: begin
        IMAGE_addr <= 5690;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5550;
        test_state <= test_b1_S5707;
      end
      test_b1_S5707: begin
        IMAGE_addr <= 5691;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S5708;
      end
      test_b1_S5708: begin
        IMAGE_addr <= 5692;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5709;
      end
      test_b1_S5709: begin
        IMAGE_addr <= 5693;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4705;
        test_state <= test_b1_S5710;
      end
      test_b1_S5710: begin
        IMAGE_addr <= 5694;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 790;
        test_state <= test_b1_S5711;
      end
      test_b1_S5711: begin
        IMAGE_addr <= 5695;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S5712;
      end
      test_b1_S5712: begin
        IMAGE_addr <= 5696;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5705;
        test_state <= test_b1_S5713;
      end
      test_b1_S5713: begin
        IMAGE_addr <= 5697;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5714;
      end
      test_b1_S5714: begin
        IMAGE_addr <= 5698;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5552;
        test_state <= test_b1_S5715;
      end
      test_b1_S5715: begin
        IMAGE_addr <= 5699;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 155;
        test_state <= test_b1_S5716;
      end
      test_b1_S5716: begin
        IMAGE_addr <= 5700;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5717;
      end
      test_b1_S5717: begin
        IMAGE_addr <= 5701;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5551;
        test_state <= test_b1_S5718;
      end
      test_b1_S5718: begin
        IMAGE_addr <= 5702;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S5719;
      end
      test_b1_S5719: begin
        IMAGE_addr <= 5703;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5605;
        test_state <= test_b1_S5720;
      end
      test_b1_S5720: begin
        IMAGE_addr <= 5704;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5721;
      end
      test_b1_S5721: begin
        IMAGE_addr <= 5705;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S5722;
      end
      test_b1_S5722: begin
        IMAGE_addr <= 5706;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5724;
        test_state <= test_b1_S5723;
      end
      test_b1_S5723: begin
        IMAGE_addr <= 5707;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5724;
      end
      test_b1_S5724: begin
        IMAGE_addr <= 5708;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5551;
        test_state <= test_b1_S5725;
      end
      test_b1_S5725: begin
        IMAGE_addr <= 5709;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S5726;
      end
      test_b1_S5726: begin
        IMAGE_addr <= 5710;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1232;
        test_state <= test_b1_S5727;
      end
      test_b1_S5727: begin
        IMAGE_addr <= 5711;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S5728;
      end
      test_b1_S5728: begin
        IMAGE_addr <= 5712;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5720;
        test_state <= test_b1_S5729;
      end
      test_b1_S5729: begin
        IMAGE_addr <= 5713;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 583;
        test_state <= test_b1_S5730;
      end
      test_b1_S5730: begin
        IMAGE_addr <= 5714;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S5731;
      end
      test_b1_S5731: begin
        IMAGE_addr <= 5715;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5605;
        test_state <= test_b1_S5732;
      end
      test_b1_S5732: begin
        IMAGE_addr <= 5716;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5733;
      end
      test_b1_S5733: begin
        IMAGE_addr <= 5717;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5552;
        test_state <= test_b1_S5734;
      end
      test_b1_S5734: begin
        IMAGE_addr <= 5718;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 155;
        test_state <= test_b1_S5735;
      end
      test_b1_S5735: begin
        IMAGE_addr <= 5719;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5736;
      end
      test_b1_S5736: begin
        IMAGE_addr <= 5720;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5737;
      end
      test_b1_S5737: begin
        IMAGE_addr <= 5721;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 52;
        test_state <= test_b1_S5738;
      end
      test_b1_S5738: begin
        IMAGE_addr <= 5722;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 732;
        test_state <= test_b1_S5739;
      end
      test_b1_S5739: begin
        IMAGE_addr <= 5723;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5740;
      end
      test_b1_S5740: begin
        IMAGE_addr <= 5724;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 732;
        test_state <= test_b1_S5741;
      end
      test_b1_S5741: begin
        IMAGE_addr <= 5725;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5742;
      end
      test_b1_S5742: begin
        IMAGE_addr <= 5726;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5743;
      end
      test_b1_S5743: begin
        IMAGE_addr <= 5727;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5679;
        test_state <= test_b1_S5744;
      end
      test_b1_S5744: begin
        IMAGE_addr <= 5728;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S5745;
      end
      test_b1_S5745: begin
        IMAGE_addr <= 5729;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5734;
        test_state <= test_b1_S5746;
      end
      test_b1_S5746: begin
        IMAGE_addr <= 5730;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S5747;
      end
      test_b1_S5747: begin
        IMAGE_addr <= 5731;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S5748;
      end
      test_b1_S5748: begin
        IMAGE_addr <= 5732;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 121;
        test_state <= test_b1_S5749;
      end
      test_b1_S5749: begin
        IMAGE_addr <= 5733;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S5750;
      end
      test_b1_S5750: begin
        IMAGE_addr <= 5734;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5751;
      end
      test_b1_S5751: begin
        IMAGE_addr <= 5735;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5552;
        test_state <= test_b1_S5752;
      end
      test_b1_S5752: begin
        IMAGE_addr <= 5736;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 147;
        test_state <= test_b1_S5753;
      end
      test_b1_S5753: begin
        IMAGE_addr <= 5737;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 400;
        test_state <= test_b1_S5754;
      end
      test_b1_S5754: begin
        IMAGE_addr <= 5738;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5624;
        test_state <= test_b1_S5755;
      end
      test_b1_S5755: begin
        IMAGE_addr <= 5739;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5648;
        test_state <= test_b1_S5756;
      end
      test_b1_S5756: begin
        IMAGE_addr <= 5740;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5757;
      end
      test_b1_S5757: begin
        IMAGE_addr <= 5741;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5689;
        test_state <= test_b1_S5758;
      end
      test_b1_S5758: begin
        IMAGE_addr <= 5742;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5759;
      end
      test_b1_S5759: begin
        IMAGE_addr <= 5743;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 52;
        test_state <= test_b1_S5760;
      end
      test_b1_S5760: begin
        IMAGE_addr <= 5744;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 732;
        test_state <= test_b1_S5761;
      end
      test_b1_S5761: begin
        IMAGE_addr <= 5745;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5762;
      end
      test_b1_S5762: begin
        IMAGE_addr <= 5746;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5552;
        test_state <= test_b1_S5763;
      end
      test_b1_S5763: begin
        IMAGE_addr <= 5747;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S5764;
      end
      test_b1_S5764: begin
        IMAGE_addr <= 5748;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5765;
      end
      test_b1_S5765: begin
        IMAGE_addr <= 5749;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5766;
      end
      test_b1_S5766: begin
        IMAGE_addr <= 5750;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5247;
        test_state <= test_b1_S5767;
      end
      test_b1_S5767: begin
        IMAGE_addr <= 5751;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S5768;
      end
      test_b1_S5768: begin
        IMAGE_addr <= 5752;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5761;
        test_state <= test_b1_S5769;
      end
      test_b1_S5769: begin
        IMAGE_addr <= 5753;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 98;
        test_state <= test_b1_S5770;
      end
      test_b1_S5770: begin
        IMAGE_addr <= 5754;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 117;
        test_state <= test_b1_S5771;
      end
      test_b1_S5771: begin
        IMAGE_addr <= 5755;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 102;
        test_state <= test_b1_S5772;
      end
      test_b1_S5772: begin
        IMAGE_addr <= 5756;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 102;
        test_state <= test_b1_S5773;
      end
      test_b1_S5773: begin
        IMAGE_addr <= 5757;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S5774;
      end
      test_b1_S5774: begin
        IMAGE_addr <= 5758;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S5775;
      end
      test_b1_S5775: begin
        IMAGE_addr <= 5759;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S5776;
      end
      test_b1_S5776: begin
        IMAGE_addr <= 5760;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S5777;
      end
      test_b1_S5777: begin
        IMAGE_addr <= 5761;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 909;
        test_state <= test_b1_S5778;
      end
      test_b1_S5778: begin
        IMAGE_addr <= 5762;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5779;
      end
      test_b1_S5779: begin
        IMAGE_addr <= 5763;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S5780;
      end
      test_b1_S5780: begin
        IMAGE_addr <= 5764;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 18;
        test_state <= test_b1_S5781;
      end
      test_b1_S5781: begin
        IMAGE_addr <= 5765;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 206;
        test_state <= test_b1_S5782;
      end
      test_b1_S5782: begin
        IMAGE_addr <= 5766;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 16;
        test_state <= test_b1_S5783;
      end
      test_b1_S5783: begin
        IMAGE_addr <= 5767;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5784;
      end
      test_b1_S5784: begin
        IMAGE_addr <= 5768;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5785;
      end
      test_b1_S5785: begin
        IMAGE_addr <= 5769;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5750;
        test_state <= test_b1_S5786;
      end
      test_b1_S5786: begin
        IMAGE_addr <= 5770;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 310;
        test_state <= test_b1_S5787;
      end
      test_b1_S5787: begin
        IMAGE_addr <= 5771;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5777;
        test_state <= test_b1_S5788;
      end
      test_b1_S5788: begin
        IMAGE_addr <= 5772;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 110;
        test_state <= test_b1_S5789;
      end
      test_b1_S5789: begin
        IMAGE_addr <= 5773;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S5790;
      end
      test_b1_S5790: begin
        IMAGE_addr <= 5774;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 120;
        test_state <= test_b1_S5791;
      end
      test_b1_S5791: begin
        IMAGE_addr <= 5775;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S5792;
      end
      test_b1_S5792: begin
        IMAGE_addr <= 5776;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S5793;
      end
      test_b1_S5793: begin
        IMAGE_addr <= 5777;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6;
        test_state <= test_b1_S5794;
      end
      test_b1_S5794: begin
        IMAGE_addr <= 5778;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5247;
        test_state <= test_b1_S5795;
      end
      test_b1_S5795: begin
        IMAGE_addr <= 5779;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S5796;
      end
      test_b1_S5796: begin
        IMAGE_addr <= 5780;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5792;
        test_state <= test_b1_S5797;
      end
      test_b1_S5797: begin
        IMAGE_addr <= 5781;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S5798;
      end
      test_b1_S5798: begin
        IMAGE_addr <= 5782;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S5799;
      end
      test_b1_S5799: begin
        IMAGE_addr <= 5783;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 109;
        test_state <= test_b1_S5800;
      end
      test_b1_S5800: begin
        IMAGE_addr <= 5784;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 112;
        test_state <= test_b1_S5801;
      end
      test_b1_S5801: begin
        IMAGE_addr <= 5785;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 83;
        test_state <= test_b1_S5802;
      end
      test_b1_S5802: begin
        IMAGE_addr <= 5786;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S5803;
      end
      test_b1_S5803: begin
        IMAGE_addr <= 5787;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S5804;
      end
      test_b1_S5804: begin
        IMAGE_addr <= 5788;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S5805;
      end
      test_b1_S5805: begin
        IMAGE_addr <= 5789;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 110;
        test_state <= test_b1_S5806;
      end
      test_b1_S5806: begin
        IMAGE_addr <= 5790;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 103;
        test_state <= test_b1_S5807;
      end
      test_b1_S5807: begin
        IMAGE_addr <= 5791;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S5808;
      end
      test_b1_S5808: begin
        IMAGE_addr <= 5792;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S5809;
      end
      test_b1_S5809: begin
        IMAGE_addr <= 5793;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S5810;
      end
      test_b1_S5810: begin
        IMAGE_addr <= 5794;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 886;
        test_state <= test_b1_S5811;
      end
      test_b1_S5811: begin
        IMAGE_addr <= 5795;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 26;
        test_state <= test_b1_S5812;
      end
      test_b1_S5812: begin
        IMAGE_addr <= 5796;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5813;
      end
      test_b1_S5813: begin
        IMAGE_addr <= 5797;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5777;
        test_state <= test_b1_S5814;
      end
      test_b1_S5814: begin
        IMAGE_addr <= 5798;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S5815;
      end
      test_b1_S5815: begin
        IMAGE_addr <= 5799;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 915;
        test_state <= test_b1_S5816;
      end
      test_b1_S5816: begin
        IMAGE_addr <= 5800;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 790;
        test_state <= test_b1_S5817;
      end
      test_b1_S5817: begin
        IMAGE_addr <= 5801;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S5818;
      end
      test_b1_S5818: begin
        IMAGE_addr <= 5802;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5809;
        test_state <= test_b1_S5819;
      end
      test_b1_S5819: begin
        IMAGE_addr <= 5803;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5820;
      end
      test_b1_S5820: begin
        IMAGE_addr <= 5804;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S5821;
      end
      test_b1_S5821: begin
        IMAGE_addr <= 5805;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5822;
      end
      test_b1_S5822: begin
        IMAGE_addr <= 5806;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5777;
        test_state <= test_b1_S5823;
      end
      test_b1_S5823: begin
        IMAGE_addr <= 5807;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S5824;
      end
      test_b1_S5824: begin
        IMAGE_addr <= 5808;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5825;
      end
      test_b1_S5825: begin
        IMAGE_addr <= 5809;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 751;
        test_state <= test_b1_S5826;
      end
      test_b1_S5826: begin
        IMAGE_addr <= 5810;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5827;
      end
      test_b1_S5827: begin
        IMAGE_addr <= 5811;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5777;
        test_state <= test_b1_S5828;
      end
      test_b1_S5828: begin
        IMAGE_addr <= 5812;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S5829;
      end
      test_b1_S5829: begin
        IMAGE_addr <= 5813;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 909;
        test_state <= test_b1_S5830;
      end
      test_b1_S5830: begin
        IMAGE_addr <= 5814;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 18;
        test_state <= test_b1_S5831;
      end
      test_b1_S5831: begin
        IMAGE_addr <= 5815;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5761;
        test_state <= test_b1_S5832;
      end
      test_b1_S5832: begin
        IMAGE_addr <= 5816;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 16;
        test_state <= test_b1_S5833;
      end
      test_b1_S5833: begin
        IMAGE_addr <= 5817;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S5834;
      end
      test_b1_S5834: begin
        IMAGE_addr <= 5818;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5822;
        test_state <= test_b1_S5835;
      end
      test_b1_S5835: begin
        IMAGE_addr <= 5819;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S5836;
      end
      test_b1_S5836: begin
        IMAGE_addr <= 5820;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4126;
        test_state <= test_b1_S5837;
      end
      test_b1_S5837: begin
        IMAGE_addr <= 5821;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5838;
      end
      test_b1_S5838: begin
        IMAGE_addr <= 5822;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 774;
        test_state <= test_b1_S5839;
      end
      test_b1_S5839: begin
        IMAGE_addr <= 5823;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5840;
      end
      test_b1_S5840: begin
        IMAGE_addr <= 5824;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5777;
        test_state <= test_b1_S5841;
      end
      test_b1_S5841: begin
        IMAGE_addr <= 5825;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2651;
        test_state <= test_b1_S5842;
      end
      test_b1_S5842: begin
        IMAGE_addr <= 5826;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5843;
      end
      test_b1_S5843: begin
        IMAGE_addr <= 5827;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5844;
      end
      test_b1_S5844: begin
        IMAGE_addr <= 5828;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5778;
        test_state <= test_b1_S5845;
      end
      test_b1_S5845: begin
        IMAGE_addr <= 5829;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 310;
        test_state <= test_b1_S5846;
      end
      test_b1_S5846: begin
        IMAGE_addr <= 5830;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5835;
        test_state <= test_b1_S5847;
      end
      test_b1_S5847: begin
        IMAGE_addr <= 5831;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S5848;
      end
      test_b1_S5848: begin
        IMAGE_addr <= 5832;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 110;
        test_state <= test_b1_S5849;
      end
      test_b1_S5849: begin
        IMAGE_addr <= 5833;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 100;
        test_state <= test_b1_S5850;
      end
      test_b1_S5850: begin
        IMAGE_addr <= 5834;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S5851;
      end
      test_b1_S5851: begin
        IMAGE_addr <= 5835;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2318;
        test_state <= test_b1_S5852;
      end
      test_b1_S5852: begin
        IMAGE_addr <= 5836;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5828;
        test_state <= test_b1_S5853;
      end
      test_b1_S5853: begin
        IMAGE_addr <= 5837;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S5854;
      end
      test_b1_S5854: begin
        IMAGE_addr <= 5838;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5843;
        test_state <= test_b1_S5855;
      end
      test_b1_S5855: begin
        IMAGE_addr <= 5839;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 112;
        test_state <= test_b1_S5856;
      end
      test_b1_S5856: begin
        IMAGE_addr <= 5840;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S5857;
      end
      test_b1_S5857: begin
        IMAGE_addr <= 5841;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 100;
        test_state <= test_b1_S5858;
      end
      test_b1_S5858: begin
        IMAGE_addr <= 5842;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S5859;
      end
      test_b1_S5859: begin
        IMAGE_addr <= 5843;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 909;
        test_state <= test_b1_S5860;
      end
      test_b1_S5860: begin
        IMAGE_addr <= 5844;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5861;
      end
      test_b1_S5861: begin
        IMAGE_addr <= 5845;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S5862;
      end
      test_b1_S5862: begin
        IMAGE_addr <= 5846;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 18;
        test_state <= test_b1_S5863;
      end
      test_b1_S5863: begin
        IMAGE_addr <= 5847;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 206;
        test_state <= test_b1_S5864;
      end
      test_b1_S5864: begin
        IMAGE_addr <= 5848;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 16;
        test_state <= test_b1_S5865;
      end
      test_b1_S5865: begin
        IMAGE_addr <= 5849;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5866;
      end
      test_b1_S5866: begin
        IMAGE_addr <= 5850;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5867;
      end
      test_b1_S5867: begin
        IMAGE_addr <= 5851;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5836;
        test_state <= test_b1_S5868;
      end
      test_b1_S5868: begin
        IMAGE_addr <= 5852;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S5869;
      end
      test_b1_S5869: begin
        IMAGE_addr <= 5853;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5859;
        test_state <= test_b1_S5870;
      end
      test_b1_S5870: begin
        IMAGE_addr <= 5854;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 107;
        test_state <= test_b1_S5871;
      end
      test_b1_S5871: begin
        IMAGE_addr <= 5855;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S5872;
      end
      test_b1_S5872: begin
        IMAGE_addr <= 5856;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S5873;
      end
      test_b1_S5873: begin
        IMAGE_addr <= 5857;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 112;
        test_state <= test_b1_S5874;
      end
      test_b1_S5874: begin
        IMAGE_addr <= 5858;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S5875;
      end
      test_b1_S5875: begin
        IMAGE_addr <= 5859;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5876;
      end
      test_b1_S5876: begin
        IMAGE_addr <= 5860;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S5877;
      end
      test_b1_S5877: begin
        IMAGE_addr <= 5861;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S5878;
      end
      test_b1_S5878: begin
        IMAGE_addr <= 5862;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5879;
      end
      test_b1_S5879: begin
        IMAGE_addr <= 5863;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 892;
        test_state <= test_b1_S5880;
      end
      test_b1_S5880: begin
        IMAGE_addr <= 5864;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5881;
      end
      test_b1_S5881: begin
        IMAGE_addr <= 5865;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5792;
        test_state <= test_b1_S5882;
      end
      test_b1_S5882: begin
        IMAGE_addr <= 5866;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 732;
        test_state <= test_b1_S5883;
      end
      test_b1_S5883: begin
        IMAGE_addr <= 5867;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 310;
        test_state <= test_b1_S5884;
      end
      test_b1_S5884: begin
        IMAGE_addr <= 5868;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5885;
      end
      test_b1_S5885: begin
        IMAGE_addr <= 5869;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5886;
      end
      test_b1_S5886: begin
        IMAGE_addr <= 5870;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5851;
        test_state <= test_b1_S5887;
      end
      test_b1_S5887: begin
        IMAGE_addr <= 5871;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S5888;
      end
      test_b1_S5888: begin
        IMAGE_addr <= 5872;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5878;
        test_state <= test_b1_S5889;
      end
      test_b1_S5889: begin
        IMAGE_addr <= 5873;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 62;
        test_state <= test_b1_S5890;
      end
      test_b1_S5890: begin
        IMAGE_addr <= 5874;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 112;
        test_state <= test_b1_S5891;
      end
      test_b1_S5891: begin
        IMAGE_addr <= 5875;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S5892;
      end
      test_b1_S5892: begin
        IMAGE_addr <= 5876;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 100;
        test_state <= test_b1_S5893;
      end
      test_b1_S5893: begin
        IMAGE_addr <= 5877;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S5894;
      end
      test_b1_S5894: begin
        IMAGE_addr <= 5878;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5843;
        test_state <= test_b1_S5895;
      end
      test_b1_S5895: begin
        IMAGE_addr <= 5879;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 132;
        test_state <= test_b1_S5896;
      end
      test_b1_S5896: begin
        IMAGE_addr <= 5880;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 877;
        test_state <= test_b1_S5897;
      end
      test_b1_S5897: begin
        IMAGE_addr <= 5881;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 26;
        test_state <= test_b1_S5898;
      end
      test_b1_S5898: begin
        IMAGE_addr <= 5882;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4126;
        test_state <= test_b1_S5899;
      end
      test_b1_S5899: begin
        IMAGE_addr <= 5883;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5843;
        test_state <= test_b1_S5900;
      end
      test_b1_S5900: begin
        IMAGE_addr <= 5884;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5859;
        test_state <= test_b1_S5901;
      end
      test_b1_S5901: begin
        IMAGE_addr <= 5885;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5902;
      end
      test_b1_S5902: begin
        IMAGE_addr <= 5886;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5903;
      end
      test_b1_S5903: begin
        IMAGE_addr <= 5887;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5870;
        test_state <= test_b1_S5904;
      end
      test_b1_S5904: begin
        IMAGE_addr <= 5888;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S5905;
      end
      test_b1_S5905: begin
        IMAGE_addr <= 5889;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5895;
        test_state <= test_b1_S5906;
      end
      test_b1_S5906: begin
        IMAGE_addr <= 5890;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 99;
        test_state <= test_b1_S5907;
      end
      test_b1_S5907: begin
        IMAGE_addr <= 5891;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 104;
        test_state <= test_b1_S5908;
      end
      test_b1_S5908: begin
        IMAGE_addr <= 5892;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 111;
        test_state <= test_b1_S5909;
      end
      test_b1_S5909: begin
        IMAGE_addr <= 5893;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 112;
        test_state <= test_b1_S5910;
      end
      test_b1_S5910: begin
        IMAGE_addr <= 5894;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S5911;
      end
      test_b1_S5911: begin
        IMAGE_addr <= 5895;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5912;
      end
      test_b1_S5912: begin
        IMAGE_addr <= 5896;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5835;
        test_state <= test_b1_S5913;
      end
      test_b1_S5913: begin
        IMAGE_addr <= 5897;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2665;
        test_state <= test_b1_S5914;
      end
      test_b1_S5914: begin
        IMAGE_addr <= 5898;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5915;
      end
      test_b1_S5915: begin
        IMAGE_addr <= 5899;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S5916;
      end
      test_b1_S5916: begin
        IMAGE_addr <= 5900;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5917;
      end
      test_b1_S5917: begin
        IMAGE_addr <= 5901;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5835;
        test_state <= test_b1_S5918;
      end
      test_b1_S5918: begin
        IMAGE_addr <= 5902;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S5919;
      end
      test_b1_S5919: begin
        IMAGE_addr <= 5903;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S5920;
      end
      test_b1_S5920: begin
        IMAGE_addr <= 5904;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5921;
      end
      test_b1_S5921: begin
        IMAGE_addr <= 5905;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5922;
      end
      test_b1_S5922: begin
        IMAGE_addr <= 5906;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5887;
        test_state <= test_b1_S5923;
      end
      test_b1_S5923: begin
        IMAGE_addr <= 5907;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S5924;
      end
      test_b1_S5924: begin
        IMAGE_addr <= 5908;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5912;
        test_state <= test_b1_S5925;
      end
      test_b1_S5925: begin
        IMAGE_addr <= 5909;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 62;
        test_state <= test_b1_S5926;
      end
      test_b1_S5926: begin
        IMAGE_addr <= 5910;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 36;
        test_state <= test_b1_S5927;
      end
      test_b1_S5927: begin
        IMAGE_addr <= 5911;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S5928;
      end
      test_b1_S5928: begin
        IMAGE_addr <= 5912;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S5929;
      end
      test_b1_S5929: begin
        IMAGE_addr <= 5913;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5930;
      end
      test_b1_S5930: begin
        IMAGE_addr <= 5914;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8;
        test_state <= test_b1_S5931;
      end
      test_b1_S5931: begin
        IMAGE_addr <= 5915;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 790;
        test_state <= test_b1_S5932;
      end
      test_b1_S5932: begin
        IMAGE_addr <= 5916;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S5933;
      end
      test_b1_S5933: begin
        IMAGE_addr <= 5917;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5921;
        test_state <= test_b1_S5934;
      end
      test_b1_S5934: begin
        IMAGE_addr <= 5918;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5895;
        test_state <= test_b1_S5935;
      end
      test_b1_S5935: begin
        IMAGE_addr <= 5919;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S5936;
      end
      test_b1_S5936: begin
        IMAGE_addr <= 5920;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5937;
      end
      test_b1_S5937: begin
        IMAGE_addr <= 5921;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S5938;
      end
      test_b1_S5938: begin
        IMAGE_addr <= 5922;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5931;
        test_state <= test_b1_S5939;
      end
      test_b1_S5939: begin
        IMAGE_addr <= 5923;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5940;
      end
      test_b1_S5940: begin
        IMAGE_addr <= 5924;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5835;
        test_state <= test_b1_S5941;
      end
      test_b1_S5941: begin
        IMAGE_addr <= 5925;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S5942;
      end
      test_b1_S5942: begin
        IMAGE_addr <= 5926;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 197;
        test_state <= test_b1_S5943;
      end
      test_b1_S5943: begin
        IMAGE_addr <= 5927;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5944;
      end
      test_b1_S5944: begin
        IMAGE_addr <= 5928;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5835;
        test_state <= test_b1_S5945;
      end
      test_b1_S5945: begin
        IMAGE_addr <= 5929;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S5946;
      end
      test_b1_S5946: begin
        IMAGE_addr <= 5930;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5947;
      end
      test_b1_S5947: begin
        IMAGE_addr <= 5931;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 732;
        test_state <= test_b1_S5948;
      end
      test_b1_S5948: begin
        IMAGE_addr <= 5932;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5949;
      end
      test_b1_S5949: begin
        IMAGE_addr <= 5933;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5950;
      end
      test_b1_S5950: begin
        IMAGE_addr <= 5934;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5906;
        test_state <= test_b1_S5951;
      end
      test_b1_S5951: begin
        IMAGE_addr <= 5935;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S5952;
      end
      test_b1_S5952: begin
        IMAGE_addr <= 5936;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5942;
        test_state <= test_b1_S5953;
      end
      test_b1_S5953: begin
        IMAGE_addr <= 5937;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S5954;
      end
      test_b1_S5954: begin
        IMAGE_addr <= 5938;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 110;
        test_state <= test_b1_S5955;
      end
      test_b1_S5955: begin
        IMAGE_addr <= 5939;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 100;
        test_state <= test_b1_S5956;
      end
      test_b1_S5956: begin
        IMAGE_addr <= 5940;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 63;
        test_state <= test_b1_S5957;
      end
      test_b1_S5957: begin
        IMAGE_addr <= 5941;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S5958;
      end
      test_b1_S5958: begin
        IMAGE_addr <= 5942;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5959;
      end
      test_b1_S5959: begin
        IMAGE_addr <= 5943;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5835;
        test_state <= test_b1_S5960;
      end
      test_b1_S5960: begin
        IMAGE_addr <= 5944;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S5961;
      end
      test_b1_S5961: begin
        IMAGE_addr <= 5945;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 27;
        test_state <= test_b1_S5962;
      end
      test_b1_S5962: begin
        IMAGE_addr <= 5946;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S5963;
      end
      test_b1_S5963: begin
        IMAGE_addr <= 5947;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5964;
      end
      test_b1_S5964: begin
        IMAGE_addr <= 5948;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 34;
        test_state <= test_b1_S5965;
      end
      test_b1_S5965: begin
        IMAGE_addr <= 5949;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 790;
        test_state <= test_b1_S5966;
      end
      test_b1_S5966: begin
        IMAGE_addr <= 5950;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S5967;
      end
      test_b1_S5967: begin
        IMAGE_addr <= 5951;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5957;
        test_state <= test_b1_S5968;
      end
      test_b1_S5968: begin
        IMAGE_addr <= 5952;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5895;
        test_state <= test_b1_S5969;
      end
      test_b1_S5969: begin
        IMAGE_addr <= 5953;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5878;
        test_state <= test_b1_S5970;
      end
      test_b1_S5970: begin
        IMAGE_addr <= 5954;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5971;
      end
      test_b1_S5971: begin
        IMAGE_addr <= 5955;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4294967295;
        test_state <= test_b1_S5972;
      end
      test_b1_S5972: begin
        IMAGE_addr <= 5956;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5973;
      end
      test_b1_S5973: begin
        IMAGE_addr <= 5957;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S5974;
      end
      test_b1_S5974: begin
        IMAGE_addr <= 5958;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5962;
        test_state <= test_b1_S5975;
      end
      test_b1_S5975: begin
        IMAGE_addr <= 5959;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5976;
      end
      test_b1_S5976: begin
        IMAGE_addr <= 5960;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S5977;
      end
      test_b1_S5977: begin
        IMAGE_addr <= 5961;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5978;
      end
      test_b1_S5978: begin
        IMAGE_addr <= 5962;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 732;
        test_state <= test_b1_S5979;
      end
      test_b1_S5979: begin
        IMAGE_addr <= 5963;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5980;
      end
      test_b1_S5980: begin
        IMAGE_addr <= 5964;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5981;
      end
      test_b1_S5981: begin
        IMAGE_addr <= 5965;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5934;
        test_state <= test_b1_S5982;
      end
      test_b1_S5982: begin
        IMAGE_addr <= 5966;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S5983;
      end
      test_b1_S5983: begin
        IMAGE_addr <= 5967;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5974;
        test_state <= test_b1_S5984;
      end
      test_b1_S5984: begin
        IMAGE_addr <= 5968;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 110;
        test_state <= test_b1_S5985;
      end
      test_b1_S5985: begin
        IMAGE_addr <= 5969;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 111;
        test_state <= test_b1_S5986;
      end
      test_b1_S5986: begin
        IMAGE_addr <= 5970;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 69;
        test_state <= test_b1_S5987;
      end
      test_b1_S5987: begin
        IMAGE_addr <= 5971;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S5988;
      end
      test_b1_S5988: begin
        IMAGE_addr <= 5972;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S5989;
      end
      test_b1_S5989: begin
        IMAGE_addr <= 5973;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S5990;
      end
      test_b1_S5990: begin
        IMAGE_addr <= 5974;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5991;
      end
      test_b1_S5991: begin
        IMAGE_addr <= 5975;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 398;
        test_state <= test_b1_S5992;
      end
      test_b1_S5992: begin
        IMAGE_addr <= 5976;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 155;
        test_state <= test_b1_S5993;
      end
      test_b1_S5993: begin
        IMAGE_addr <= 5977;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 183;
        test_state <= test_b1_S5994;
      end
      test_b1_S5994: begin
        IMAGE_addr <= 5978;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S5995;
      end
      test_b1_S5995: begin
        IMAGE_addr <= 5979;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 398;
        test_state <= test_b1_S5996;
      end
      test_b1_S5996: begin
        IMAGE_addr <= 5980;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 147;
        test_state <= test_b1_S5997;
      end
      test_b1_S5997: begin
        IMAGE_addr <= 5981;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5998;
      end
      test_b1_S5998: begin
        IMAGE_addr <= 5982;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S5999;
      end
      test_b1_S5999: begin
        IMAGE_addr <= 5983;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5965;
        test_state <= test_b1_S6000;
      end
      test_b1_S6000: begin
        IMAGE_addr <= 5984;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S6001;
      end
      test_b1_S6001: begin
        IMAGE_addr <= 5985;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5994;
        test_state <= test_b1_S6002;
      end
      test_b1_S6002: begin
        IMAGE_addr <= 5986;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 119;
        test_state <= test_b1_S6003;
      end
      test_b1_S6003: begin
        IMAGE_addr <= 5987;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S6004;
      end
      test_b1_S6004: begin
        IMAGE_addr <= 5988;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S6005;
      end
      test_b1_S6005: begin
        IMAGE_addr <= 5989;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 104;
        test_state <= test_b1_S6006;
      end
      test_b1_S6006: begin
        IMAGE_addr <= 5990;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 80;
        test_state <= test_b1_S6007;
      end
      test_b1_S6007: begin
        IMAGE_addr <= 5991;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S6008;
      end
      test_b1_S6008: begin
        IMAGE_addr <= 5992;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 100;
        test_state <= test_b1_S6009;
      end
      test_b1_S6009: begin
        IMAGE_addr <= 5993;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6010;
      end
      test_b1_S6010: begin
        IMAGE_addr <= 5994;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6011;
      end
      test_b1_S6011: begin
        IMAGE_addr <= 5995;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 32;
        test_state <= test_b1_S6012;
      end
      test_b1_S6012: begin
        IMAGE_addr <= 5996;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5843;
        test_state <= test_b1_S6013;
      end
      test_b1_S6013: begin
        IMAGE_addr <= 5997;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 27;
        test_state <= test_b1_S6014;
      end
      test_b1_S6014: begin
        IMAGE_addr <= 5998;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S6015;
      end
      test_b1_S6015: begin
        IMAGE_addr <= 5999;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6016;
      end
      test_b1_S6016: begin
        IMAGE_addr <= 6000;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5843;
        test_state <= test_b1_S6017;
      end
      test_b1_S6017: begin
        IMAGE_addr <= 6001;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6018;
      end
      test_b1_S6018: begin
        IMAGE_addr <= 6002;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 400;
        test_state <= test_b1_S6019;
      end
      test_b1_S6019: begin
        IMAGE_addr <= 6003;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2820;
        test_state <= test_b1_S6020;
      end
      test_b1_S6020: begin
        IMAGE_addr <= 6004;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5974;
        test_state <= test_b1_S6021;
      end
      test_b1_S6021: begin
        IMAGE_addr <= 6005;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6022;
      end
      test_b1_S6022: begin
        IMAGE_addr <= 6006;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 400;
        test_state <= test_b1_S6023;
      end
      test_b1_S6023: begin
        IMAGE_addr <= 6007;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2801;
        test_state <= test_b1_S6024;
      end
      test_b1_S6024: begin
        IMAGE_addr <= 6008;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6025;
      end
      test_b1_S6025: begin
        IMAGE_addr <= 6009;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6026;
      end
      test_b1_S6026: begin
        IMAGE_addr <= 6010;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5983;
        test_state <= test_b1_S6027;
      end
      test_b1_S6027: begin
        IMAGE_addr <= 6011;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S6028;
      end
      test_b1_S6028: begin
        IMAGE_addr <= 6012;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6017;
        test_state <= test_b1_S6029;
      end
      test_b1_S6029: begin
        IMAGE_addr <= 6013;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 103;
        test_state <= test_b1_S6030;
      end
      test_b1_S6030: begin
        IMAGE_addr <= 6014;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S6031;
      end
      test_b1_S6031: begin
        IMAGE_addr <= 6015;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S6032;
      end
      test_b1_S6032: begin
        IMAGE_addr <= 6016;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6033;
      end
      test_b1_S6033: begin
        IMAGE_addr <= 6017;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 466;
        test_state <= test_b1_S6034;
      end
      test_b1_S6034: begin
        IMAGE_addr <= 6018;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S6035;
      end
      test_b1_S6035: begin
        IMAGE_addr <= 6019;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 359;
        test_state <= test_b1_S6036;
      end
      test_b1_S6036: begin
        IMAGE_addr <= 6020;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6037;
      end
      test_b1_S6037: begin
        IMAGE_addr <= 6021;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6038;
      end
      test_b1_S6038: begin
        IMAGE_addr <= 6022;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5778;
        test_state <= test_b1_S6039;
      end
      test_b1_S6039: begin
        IMAGE_addr <= 6023;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4705;
        test_state <= test_b1_S6040;
      end
      test_b1_S6040: begin
        IMAGE_addr <= 6024;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6029;
        test_state <= test_b1_S6041;
      end
      test_b1_S6041: begin
        IMAGE_addr <= 6025;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 95;
        test_state <= test_b1_S6042;
      end
      test_b1_S6042: begin
        IMAGE_addr <= 6026;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 95;
        test_state <= test_b1_S6043;
      end
      test_b1_S6043: begin
        IMAGE_addr <= 6027;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 34;
        test_state <= test_b1_S6044;
      end
      test_b1_S6044: begin
        IMAGE_addr <= 6028;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6045;
      end
      test_b1_S6045: begin
        IMAGE_addr <= 6029;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6046;
      end
      test_b1_S6046: begin
        IMAGE_addr <= 6030;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6047;
      end
      test_b1_S6047: begin
        IMAGE_addr <= 6031;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S6048;
      end
      test_b1_S6048: begin
        IMAGE_addr <= 6032;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 886;
        test_state <= test_b1_S6049;
      end
      test_b1_S6049: begin
        IMAGE_addr <= 6033;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 16;
        test_state <= test_b1_S6050;
      end
      test_b1_S6050: begin
        IMAGE_addr <= 6034;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6051;
      end
      test_b1_S6051: begin
        IMAGE_addr <= 6035;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5835;
        test_state <= test_b1_S6052;
      end
      test_b1_S6052: begin
        IMAGE_addr <= 6036;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S6053;
      end
      test_b1_S6053: begin
        IMAGE_addr <= 6037;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5942;
        test_state <= test_b1_S6054;
      end
      test_b1_S6054: begin
        IMAGE_addr <= 6038;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S6055;
      end
      test_b1_S6055: begin
        IMAGE_addr <= 6039;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6062;
        test_state <= test_b1_S6056;
      end
      test_b1_S6056: begin
        IMAGE_addr <= 6040;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6057;
      end
      test_b1_S6057: begin
        IMAGE_addr <= 6041;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 32;
        test_state <= test_b1_S6058;
      end
      test_b1_S6058: begin
        IMAGE_addr <= 6042;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5912;
        test_state <= test_b1_S6059;
      end
      test_b1_S6059: begin
        IMAGE_addr <= 6043;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S6060;
      end
      test_b1_S6060: begin
        IMAGE_addr <= 6044;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6060;
        test_state <= test_b1_S6061;
      end
      test_b1_S6061: begin
        IMAGE_addr <= 6045;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5942;
        test_state <= test_b1_S6062;
      end
      test_b1_S6062: begin
        IMAGE_addr <= 6046;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S6063;
      end
      test_b1_S6063: begin
        IMAGE_addr <= 6047;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6051;
        test_state <= test_b1_S6064;
      end
      test_b1_S6064: begin
        IMAGE_addr <= 6048;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6065;
      end
      test_b1_S6065: begin
        IMAGE_addr <= 6049;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6066;
      end
      test_b1_S6066: begin
        IMAGE_addr <= 6050;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6067;
      end
      test_b1_S6067: begin
        IMAGE_addr <= 6051;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S6068;
      end
      test_b1_S6068: begin
        IMAGE_addr <= 6052;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6058;
        test_state <= test_b1_S6069;
      end
      test_b1_S6069: begin
        IMAGE_addr <= 6053;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6017;
        test_state <= test_b1_S6070;
      end
      test_b1_S6070: begin
        IMAGE_addr <= 6054;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5912;
        test_state <= test_b1_S6071;
      end
      test_b1_S6071: begin
        IMAGE_addr <= 6055;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6072;
      end
      test_b1_S6072: begin
        IMAGE_addr <= 6056;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4294967295;
        test_state <= test_b1_S6073;
      end
      test_b1_S6073: begin
        IMAGE_addr <= 6057;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6074;
      end
      test_b1_S6074: begin
        IMAGE_addr <= 6058;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 732;
        test_state <= test_b1_S6075;
      end
      test_b1_S6075: begin
        IMAGE_addr <= 6059;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6076;
      end
      test_b1_S6076: begin
        IMAGE_addr <= 6060;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3433;
        test_state <= test_b1_S6077;
      end
      test_b1_S6077: begin
        IMAGE_addr <= 6061;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6078;
      end
      test_b1_S6078: begin
        IMAGE_addr <= 6062;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 758;
        test_state <= test_b1_S6079;
      end
      test_b1_S6079: begin
        IMAGE_addr <= 6063;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6080;
      end
      test_b1_S6080: begin
        IMAGE_addr <= 6064;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6081;
      end
      test_b1_S6081: begin
        IMAGE_addr <= 6065;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6022;
        test_state <= test_b1_S6082;
      end
      test_b1_S6082: begin
        IMAGE_addr <= 6066;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 306;
        test_state <= test_b1_S6083;
      end
      test_b1_S6083: begin
        IMAGE_addr <= 6067;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6070;
        test_state <= test_b1_S6084;
      end
      test_b1_S6084: begin
        IMAGE_addr <= 6068;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 34;
        test_state <= test_b1_S6085;
      end
      test_b1_S6085: begin
        IMAGE_addr <= 6069;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6086;
      end
      test_b1_S6086: begin
        IMAGE_addr <= 6070;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6087;
      end
      test_b1_S6087: begin
        IMAGE_addr <= 6071;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6088;
      end
      test_b1_S6088: begin
        IMAGE_addr <= 6072;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S6089;
      end
      test_b1_S6089: begin
        IMAGE_addr <= 6073;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6081;
        test_state <= test_b1_S6090;
      end
      test_b1_S6090: begin
        IMAGE_addr <= 6074;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6091;
      end
      test_b1_S6091: begin
        IMAGE_addr <= 6075;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 34;
        test_state <= test_b1_S6092;
      end
      test_b1_S6092: begin
        IMAGE_addr <= 6076;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 562;
        test_state <= test_b1_S6093;
      end
      test_b1_S6093: begin
        IMAGE_addr <= 6077;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5843;
        test_state <= test_b1_S6094;
      end
      test_b1_S6094: begin
        IMAGE_addr <= 6078;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 27;
        test_state <= test_b1_S6095;
      end
      test_b1_S6095: begin
        IMAGE_addr <= 6079;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5859;
        test_state <= test_b1_S6096;
      end
      test_b1_S6096: begin
        IMAGE_addr <= 6080;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6097;
      end
      test_b1_S6097: begin
        IMAGE_addr <= 6081;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5994;
        test_state <= test_b1_S6098;
      end
      test_b1_S6098: begin
        IMAGE_addr <= 6082;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6099;
      end
      test_b1_S6099: begin
        IMAGE_addr <= 6083;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6100;
      end
      test_b1_S6100: begin
        IMAGE_addr <= 6084;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6065;
        test_state <= test_b1_S6101;
      end
      test_b1_S6101: begin
        IMAGE_addr <= 6085;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 310;
        test_state <= test_b1_S6102;
      end
      test_b1_S6102: begin
        IMAGE_addr <= 6086;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6097;
        test_state <= test_b1_S6103;
      end
      test_b1_S6103: begin
        IMAGE_addr <= 6087;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 102;
        test_state <= test_b1_S6104;
      end
      test_b1_S6104: begin
        IMAGE_addr <= 6088;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 111;
        test_state <= test_b1_S6105;
      end
      test_b1_S6105: begin
        IMAGE_addr <= 6089;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S6106;
      end
      test_b1_S6106: begin
        IMAGE_addr <= 6090;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 109;
        test_state <= test_b1_S6107;
      end
      test_b1_S6107: begin
        IMAGE_addr <= 6091;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S6108;
      end
      test_b1_S6108: begin
        IMAGE_addr <= 6092;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S6109;
      end
      test_b1_S6109: begin
        IMAGE_addr <= 6093;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S6110;
      end
      test_b1_S6110: begin
        IMAGE_addr <= 6094;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S6111;
      end
      test_b1_S6111: begin
        IMAGE_addr <= 6095;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 100;
        test_state <= test_b1_S6112;
      end
      test_b1_S6112: begin
        IMAGE_addr <= 6096;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6113;
      end
      test_b1_S6113: begin
        IMAGE_addr <= 6097;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4294967295;
        test_state <= test_b1_S6114;
      end
      test_b1_S6114: begin
        IMAGE_addr <= 6098;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6084;
        test_state <= test_b1_S6115;
      end
      test_b1_S6115: begin
        IMAGE_addr <= 6099;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S6116;
      end
      test_b1_S6116: begin
        IMAGE_addr <= 6100;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6110;
        test_state <= test_b1_S6117;
      end
      test_b1_S6117: begin
        IMAGE_addr <= 6101;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 119;
        test_state <= test_b1_S6118;
      end
      test_b1_S6118: begin
        IMAGE_addr <= 6102;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S6119;
      end
      test_b1_S6119: begin
        IMAGE_addr <= 6103;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S6120;
      end
      test_b1_S6120: begin
        IMAGE_addr <= 6104;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 104;
        test_state <= test_b1_S6121;
      end
      test_b1_S6121: begin
        IMAGE_addr <= 6105;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 66;
        test_state <= test_b1_S6122;
      end
      test_b1_S6122: begin
        IMAGE_addr <= 6106;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S6123;
      end
      test_b1_S6123: begin
        IMAGE_addr <= 6107;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S6124;
      end
      test_b1_S6124: begin
        IMAGE_addr <= 6108;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S6125;
      end
      test_b1_S6125: begin
        IMAGE_addr <= 6109;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6126;
      end
      test_b1_S6126: begin
        IMAGE_addr <= 6110;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6127;
      end
      test_b1_S6127: begin
        IMAGE_addr <= 6111;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 47;
        test_state <= test_b1_S6128;
      end
      test_b1_S6128: begin
        IMAGE_addr <= 6112;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 766;
        test_state <= test_b1_S6129;
      end
      test_b1_S6129: begin
        IMAGE_addr <= 6113;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6130;
      end
      test_b1_S6130: begin
        IMAGE_addr <= 6114;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 925;
        test_state <= test_b1_S6131;
      end
      test_b1_S6131: begin
        IMAGE_addr <= 6115;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6132;
      end
      test_b1_S6132: begin
        IMAGE_addr <= 6116;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 183;
        test_state <= test_b1_S6133;
      end
      test_b1_S6133: begin
        IMAGE_addr <= 6117;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3673;
        test_state <= test_b1_S6134;
      end
      test_b1_S6134: begin
        IMAGE_addr <= 6118;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6135;
      end
      test_b1_S6135: begin
        IMAGE_addr <= 6119;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6136;
      end
      test_b1_S6136: begin
        IMAGE_addr <= 6120;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6098;
        test_state <= test_b1_S6137;
      end
      test_b1_S6137: begin
        IMAGE_addr <= 6121;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S6138;
      end
      test_b1_S6138: begin
        IMAGE_addr <= 6122;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6128;
        test_state <= test_b1_S6139;
      end
      test_b1_S6139: begin
        IMAGE_addr <= 6123;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 99;
        test_state <= test_b1_S6140;
      end
      test_b1_S6140: begin
        IMAGE_addr <= 6124;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 104;
        test_state <= test_b1_S6141;
      end
      test_b1_S6141: begin
        IMAGE_addr <= 6125;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S6142;
      end
      test_b1_S6142: begin
        IMAGE_addr <= 6126;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S6143;
      end
      test_b1_S6143: begin
        IMAGE_addr <= 6127;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6144;
      end
      test_b1_S6144: begin
        IMAGE_addr <= 6128;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 189;
        test_state <= test_b1_S6145;
      end
      test_b1_S6145: begin
        IMAGE_addr <= 6129;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S6146;
      end
      test_b1_S6146: begin
        IMAGE_addr <= 6130;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6135;
        test_state <= test_b1_S6147;
      end
      test_b1_S6147: begin
        IMAGE_addr <= 6131;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6148;
      end
      test_b1_S6148: begin
        IMAGE_addr <= 6132;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 110;
        test_state <= test_b1_S6149;
      end
      test_b1_S6149: begin
        IMAGE_addr <= 6133;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 790;
        test_state <= test_b1_S6150;
      end
      test_b1_S6150: begin
        IMAGE_addr <= 6134;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6151;
      end
      test_b1_S6151: begin
        IMAGE_addr <= 6135;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S6152;
      end
      test_b1_S6152: begin
        IMAGE_addr <= 6136;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6139;
        test_state <= test_b1_S6153;
      end
      test_b1_S6153: begin
        IMAGE_addr <= 6137;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 371;
        test_state <= test_b1_S6154;
      end
      test_b1_S6154: begin
        IMAGE_addr <= 6138;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6155;
      end
      test_b1_S6155: begin
        IMAGE_addr <= 6139;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3735;
        test_state <= test_b1_S6156;
      end
      test_b1_S6156: begin
        IMAGE_addr <= 6140;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S6157;
      end
      test_b1_S6157: begin
        IMAGE_addr <= 6141;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6146;
        test_state <= test_b1_S6158;
      end
      test_b1_S6158: begin
        IMAGE_addr <= 6142;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6159;
      end
      test_b1_S6159: begin
        IMAGE_addr <= 6143;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 39;
        test_state <= test_b1_S6160;
      end
      test_b1_S6160: begin
        IMAGE_addr <= 6144;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 790;
        test_state <= test_b1_S6161;
      end
      test_b1_S6161: begin
        IMAGE_addr <= 6145;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6162;
      end
      test_b1_S6162: begin
        IMAGE_addr <= 6146;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S6163;
      end
      test_b1_S6163: begin
        IMAGE_addr <= 6147;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6152;
        test_state <= test_b1_S6164;
      end
      test_b1_S6164: begin
        IMAGE_addr <= 6148;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6165;
      end
      test_b1_S6165: begin
        IMAGE_addr <= 6149;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 34;
        test_state <= test_b1_S6166;
      end
      test_b1_S6166: begin
        IMAGE_addr <= 6150;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 359;
        test_state <= test_b1_S6167;
      end
      test_b1_S6167: begin
        IMAGE_addr <= 6151;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6168;
      end
      test_b1_S6168: begin
        IMAGE_addr <= 6152;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3735;
        test_state <= test_b1_S6169;
      end
      test_b1_S6169: begin
        IMAGE_addr <= 6153;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S6170;
      end
      test_b1_S6170: begin
        IMAGE_addr <= 6154;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6159;
        test_state <= test_b1_S6171;
      end
      test_b1_S6171: begin
        IMAGE_addr <= 6155;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6172;
      end
      test_b1_S6172: begin
        IMAGE_addr <= 6156;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 91;
        test_state <= test_b1_S6173;
      end
      test_b1_S6173: begin
        IMAGE_addr <= 6157;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 790;
        test_state <= test_b1_S6174;
      end
      test_b1_S6174: begin
        IMAGE_addr <= 6158;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6175;
      end
      test_b1_S6175: begin
        IMAGE_addr <= 6159;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S6176;
      end
      test_b1_S6176: begin
        IMAGE_addr <= 6160;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6166;
        test_state <= test_b1_S6177;
      end
      test_b1_S6177: begin
        IMAGE_addr <= 6161;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6178;
      end
      test_b1_S6178: begin
        IMAGE_addr <= 6162;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 27;
        test_state <= test_b1_S6179;
      end
      test_b1_S6179: begin
        IMAGE_addr <= 6163;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 359;
        test_state <= test_b1_S6180;
      end
      test_b1_S6180: begin
        IMAGE_addr <= 6164;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 359;
        test_state <= test_b1_S6181;
      end
      test_b1_S6181: begin
        IMAGE_addr <= 6165;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6182;
      end
      test_b1_S6182: begin
        IMAGE_addr <= 6166;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3697;
        test_state <= test_b1_S6183;
      end
      test_b1_S6183: begin
        IMAGE_addr <= 6167;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 359;
        test_state <= test_b1_S6184;
      end
      test_b1_S6184: begin
        IMAGE_addr <= 6168;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6185;
      end
      test_b1_S6185: begin
        IMAGE_addr <= 6169;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6186;
      end
      test_b1_S6186: begin
        IMAGE_addr <= 6170;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6120;
        test_state <= test_b1_S6187;
      end
      test_b1_S6187: begin
        IMAGE_addr <= 6171;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S6188;
      end
      test_b1_S6188: begin
        IMAGE_addr <= 6172;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6177;
        test_state <= test_b1_S6189;
      end
      test_b1_S6189: begin
        IMAGE_addr <= 6173;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 111;
        test_state <= test_b1_S6190;
      end
      test_b1_S6190: begin
        IMAGE_addr <= 6174;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 98;
        test_state <= test_b1_S6191;
      end
      test_b1_S6191: begin
        IMAGE_addr <= 6175;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 106;
        test_state <= test_b1_S6192;
      end
      test_b1_S6192: begin
        IMAGE_addr <= 6176;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6193;
      end
      test_b1_S6193: begin
        IMAGE_addr <= 6177;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 189;
        test_state <= test_b1_S6194;
      end
      test_b1_S6194: begin
        IMAGE_addr <= 6178;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S6195;
      end
      test_b1_S6195: begin
        IMAGE_addr <= 6179;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6184;
        test_state <= test_b1_S6196;
      end
      test_b1_S6196: begin
        IMAGE_addr <= 6180;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6197;
      end
      test_b1_S6197: begin
        IMAGE_addr <= 6181;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 100;
        test_state <= test_b1_S6198;
      end
      test_b1_S6198: begin
        IMAGE_addr <= 6182;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 790;
        test_state <= test_b1_S6199;
      end
      test_b1_S6199: begin
        IMAGE_addr <= 6183;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6200;
      end
      test_b1_S6200: begin
        IMAGE_addr <= 6184;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S6201;
      end
      test_b1_S6201: begin
        IMAGE_addr <= 6185;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6193;
        test_state <= test_b1_S6202;
      end
      test_b1_S6202: begin
        IMAGE_addr <= 6186;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S6203;
      end
      test_b1_S6203: begin
        IMAGE_addr <= 6187;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6191;
        test_state <= test_b1_S6204;
      end
      test_b1_S6204: begin
        IMAGE_addr <= 6188;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4404;
        test_state <= test_b1_S6205;
      end
      test_b1_S6205: begin
        IMAGE_addr <= 6189;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4689;
        test_state <= test_b1_S6206;
      end
      test_b1_S6206: begin
        IMAGE_addr <= 6190;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6207;
      end
      test_b1_S6207: begin
        IMAGE_addr <= 6191;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6110;
        test_state <= test_b1_S6208;
      end
      test_b1_S6208: begin
        IMAGE_addr <= 6192;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6209;
      end
      test_b1_S6209: begin
        IMAGE_addr <= 6193;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3735;
        test_state <= test_b1_S6210;
      end
      test_b1_S6210: begin
        IMAGE_addr <= 6194;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S6211;
      end
      test_b1_S6211: begin
        IMAGE_addr <= 6195;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6200;
        test_state <= test_b1_S6212;
      end
      test_b1_S6212: begin
        IMAGE_addr <= 6196;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6213;
      end
      test_b1_S6213: begin
        IMAGE_addr <= 6197;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 111;
        test_state <= test_b1_S6214;
      end
      test_b1_S6214: begin
        IMAGE_addr <= 6198;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 790;
        test_state <= test_b1_S6215;
      end
      test_b1_S6215: begin
        IMAGE_addr <= 6199;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6216;
      end
      test_b1_S6216: begin
        IMAGE_addr <= 6200;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S6217;
      end
      test_b1_S6217: begin
        IMAGE_addr <= 6201;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6209;
        test_state <= test_b1_S6218;
      end
      test_b1_S6218: begin
        IMAGE_addr <= 6202;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S6219;
      end
      test_b1_S6219: begin
        IMAGE_addr <= 6203;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6207;
        test_state <= test_b1_S6220;
      end
      test_b1_S6220: begin
        IMAGE_addr <= 6204;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4438;
        test_state <= test_b1_S6221;
      end
      test_b1_S6221: begin
        IMAGE_addr <= 6205;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4689;
        test_state <= test_b1_S6222;
      end
      test_b1_S6222: begin
        IMAGE_addr <= 6206;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6223;
      end
      test_b1_S6223: begin
        IMAGE_addr <= 6207;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6110;
        test_state <= test_b1_S6224;
      end
      test_b1_S6224: begin
        IMAGE_addr <= 6208;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6225;
      end
      test_b1_S6225: begin
        IMAGE_addr <= 6209;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3735;
        test_state <= test_b1_S6226;
      end
      test_b1_S6226: begin
        IMAGE_addr <= 6210;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S6227;
      end
      test_b1_S6227: begin
        IMAGE_addr <= 6211;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6216;
        test_state <= test_b1_S6228;
      end
      test_b1_S6228: begin
        IMAGE_addr <= 6212;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6229;
      end
      test_b1_S6229: begin
        IMAGE_addr <= 6213;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 120;
        test_state <= test_b1_S6230;
      end
      test_b1_S6230: begin
        IMAGE_addr <= 6214;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 790;
        test_state <= test_b1_S6231;
      end
      test_b1_S6231: begin
        IMAGE_addr <= 6215;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6232;
      end
      test_b1_S6232: begin
        IMAGE_addr <= 6216;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S6233;
      end
      test_b1_S6233: begin
        IMAGE_addr <= 6217;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6225;
        test_state <= test_b1_S6234;
      end
      test_b1_S6234: begin
        IMAGE_addr <= 6218;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S6235;
      end
      test_b1_S6235: begin
        IMAGE_addr <= 6219;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6223;
        test_state <= test_b1_S6236;
      end
      test_b1_S6236: begin
        IMAGE_addr <= 6220;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4420;
        test_state <= test_b1_S6237;
      end
      test_b1_S6237: begin
        IMAGE_addr <= 6221;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4689;
        test_state <= test_b1_S6238;
      end
      test_b1_S6238: begin
        IMAGE_addr <= 6222;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6239;
      end
      test_b1_S6239: begin
        IMAGE_addr <= 6223;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6110;
        test_state <= test_b1_S6240;
      end
      test_b1_S6240: begin
        IMAGE_addr <= 6224;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6241;
      end
      test_b1_S6241: begin
        IMAGE_addr <= 6225;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3735;
        test_state <= test_b1_S6242;
      end
      test_b1_S6242: begin
        IMAGE_addr <= 6226;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S6243;
      end
      test_b1_S6243: begin
        IMAGE_addr <= 6227;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6232;
        test_state <= test_b1_S6244;
      end
      test_b1_S6244: begin
        IMAGE_addr <= 6228;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6245;
      end
      test_b1_S6245: begin
        IMAGE_addr <= 6229;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 99;
        test_state <= test_b1_S6246;
      end
      test_b1_S6246: begin
        IMAGE_addr <= 6230;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 790;
        test_state <= test_b1_S6247;
      end
      test_b1_S6247: begin
        IMAGE_addr <= 6231;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6248;
      end
      test_b1_S6248: begin
        IMAGE_addr <= 6232;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S6249;
      end
      test_b1_S6249: begin
        IMAGE_addr <= 6233;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6237;
        test_state <= test_b1_S6250;
      end
      test_b1_S6250: begin
        IMAGE_addr <= 6234;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S6251;
      end
      test_b1_S6251: begin
        IMAGE_addr <= 6235;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 359;
        test_state <= test_b1_S6252;
      end
      test_b1_S6252: begin
        IMAGE_addr <= 6236;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6253;
      end
      test_b1_S6253: begin
        IMAGE_addr <= 6237;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3735;
        test_state <= test_b1_S6254;
      end
      test_b1_S6254: begin
        IMAGE_addr <= 6238;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S6255;
      end
      test_b1_S6255: begin
        IMAGE_addr <= 6239;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6244;
        test_state <= test_b1_S6256;
      end
      test_b1_S6256: begin
        IMAGE_addr <= 6240;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6257;
      end
      test_b1_S6257: begin
        IMAGE_addr <= 6241;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S6258;
      end
      test_b1_S6258: begin
        IMAGE_addr <= 6242;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 790;
        test_state <= test_b1_S6259;
      end
      test_b1_S6259: begin
        IMAGE_addr <= 6243;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6260;
      end
      test_b1_S6260: begin
        IMAGE_addr <= 6244;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S6261;
      end
      test_b1_S6261: begin
        IMAGE_addr <= 6245;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6256;
        test_state <= test_b1_S6262;
      end
      test_b1_S6262: begin
        IMAGE_addr <= 6246;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6263;
      end
      test_b1_S6263: begin
        IMAGE_addr <= 6247;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6097;
        test_state <= test_b1_S6264;
      end
      test_b1_S6264: begin
        IMAGE_addr <= 6248;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 155;
        test_state <= test_b1_S6265;
      end
      test_b1_S6265: begin
        IMAGE_addr <= 6249;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6266;
      end
      test_b1_S6266: begin
        IMAGE_addr <= 6250;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 391;
        test_state <= test_b1_S6267;
      end
      test_b1_S6267: begin
        IMAGE_addr <= 6251;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 766;
        test_state <= test_b1_S6268;
      end
      test_b1_S6268: begin
        IMAGE_addr <= 6252;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6269;
      end
      test_b1_S6269: begin
        IMAGE_addr <= 6253;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6097;
        test_state <= test_b1_S6270;
      end
      test_b1_S6270: begin
        IMAGE_addr <= 6254;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 147;
        test_state <= test_b1_S6271;
      end
      test_b1_S6271: begin
        IMAGE_addr <= 6255;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6272;
      end
      test_b1_S6272: begin
        IMAGE_addr <= 6256;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3735;
        test_state <= test_b1_S6273;
      end
      test_b1_S6273: begin
        IMAGE_addr <= 6257;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 359;
        test_state <= test_b1_S6274;
      end
      test_b1_S6274: begin
        IMAGE_addr <= 6258;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6275;
      end
      test_b1_S6275: begin
        IMAGE_addr <= 6259;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6276;
      end
      test_b1_S6276: begin
        IMAGE_addr <= 6260;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6170;
        test_state <= test_b1_S6277;
      end
      test_b1_S6277: begin
        IMAGE_addr <= 6261;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S6278;
      end
      test_b1_S6278: begin
        IMAGE_addr <= 6262;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6271;
        test_state <= test_b1_S6279;
      end
      test_b1_S6279: begin
        IMAGE_addr <= 6263;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 99;
        test_state <= test_b1_S6280;
      end
      test_b1_S6280: begin
        IMAGE_addr <= 6264;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 111;
        test_state <= test_b1_S6281;
      end
      test_b1_S6281: begin
        IMAGE_addr <= 6265;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 109;
        test_state <= test_b1_S6282;
      end
      test_b1_S6282: begin
        IMAGE_addr <= 6266;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 112;
        test_state <= test_b1_S6283;
      end
      test_b1_S6283: begin
        IMAGE_addr <= 6267;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 108;
        test_state <= test_b1_S6284;
      end
      test_b1_S6284: begin
        IMAGE_addr <= 6268;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S6285;
      end
      test_b1_S6285: begin
        IMAGE_addr <= 6269;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 120;
        test_state <= test_b1_S6286;
      end
      test_b1_S6286: begin
        IMAGE_addr <= 6270;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6287;
      end
      test_b1_S6287: begin
        IMAGE_addr <= 6271;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 189;
        test_state <= test_b1_S6288;
      end
      test_b1_S6288: begin
        IMAGE_addr <= 6272;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 25;
        test_state <= test_b1_S6289;
      end
      test_b1_S6289: begin
        IMAGE_addr <= 6273;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S6290;
      end
      test_b1_S6290: begin
        IMAGE_addr <= 6274;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6291;
      end
      test_b1_S6291: begin
        IMAGE_addr <= 6275;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 92;
        test_state <= test_b1_S6292;
      end
      test_b1_S6292: begin
        IMAGE_addr <= 6276;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 790;
        test_state <= test_b1_S6293;
      end
      test_b1_S6293: begin
        IMAGE_addr <= 6277;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S6294;
      end
      test_b1_S6294: begin
        IMAGE_addr <= 6278;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6284;
        test_state <= test_b1_S6295;
      end
      test_b1_S6295: begin
        IMAGE_addr <= 6279;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S6296;
      end
      test_b1_S6296: begin
        IMAGE_addr <= 6280;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6128;
        test_state <= test_b1_S6297;
      end
      test_b1_S6297: begin
        IMAGE_addr <= 6281;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6298;
      end
      test_b1_S6298: begin
        IMAGE_addr <= 6282;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6299;
      end
      test_b1_S6299: begin
        IMAGE_addr <= 6283;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6300;
      end
      test_b1_S6300: begin
        IMAGE_addr <= 6284;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 751;
        test_state <= test_b1_S6301;
      end
      test_b1_S6301: begin
        IMAGE_addr <= 6285;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S6302;
      end
      test_b1_S6302: begin
        IMAGE_addr <= 6286;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6303;
      end
      test_b1_S6303: begin
        IMAGE_addr <= 6287;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 37;
        test_state <= test_b1_S6304;
      end
      test_b1_S6304: begin
        IMAGE_addr <= 6288;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 790;
        test_state <= test_b1_S6305;
      end
      test_b1_S6305: begin
        IMAGE_addr <= 6289;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S6306;
      end
      test_b1_S6306: begin
        IMAGE_addr <= 6290;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6296;
        test_state <= test_b1_S6307;
      end
      test_b1_S6307: begin
        IMAGE_addr <= 6291;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S6308;
      end
      test_b1_S6308: begin
        IMAGE_addr <= 6292;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6177;
        test_state <= test_b1_S6309;
      end
      test_b1_S6309: begin
        IMAGE_addr <= 6293;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6310;
      end
      test_b1_S6310: begin
        IMAGE_addr <= 6294;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6311;
      end
      test_b1_S6311: begin
        IMAGE_addr <= 6295;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6312;
      end
      test_b1_S6312: begin
        IMAGE_addr <= 6296;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 751;
        test_state <= test_b1_S6313;
      end
      test_b1_S6313: begin
        IMAGE_addr <= 6297;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 359;
        test_state <= test_b1_S6314;
      end
      test_b1_S6314: begin
        IMAGE_addr <= 6298;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8;
        test_state <= test_b1_S6315;
      end
      test_b1_S6315: begin
        IMAGE_addr <= 6299;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6271;
        test_state <= test_b1_S6316;
      end
      test_b1_S6316: begin
        IMAGE_addr <= 6300;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6317;
      end
      test_b1_S6317: begin
        IMAGE_addr <= 6301;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6318;
      end
      test_b1_S6318: begin
        IMAGE_addr <= 6302;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6260;
        test_state <= test_b1_S6319;
      end
      test_b1_S6319: begin
        IMAGE_addr <= 6303;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S6320;
      end
      test_b1_S6320: begin
        IMAGE_addr <= 6304;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6312;
        test_state <= test_b1_S6321;
      end
      test_b1_S6321: begin
        IMAGE_addr <= 6305;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S6322;
      end
      test_b1_S6322: begin
        IMAGE_addr <= 6306;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S6323;
      end
      test_b1_S6323: begin
        IMAGE_addr <= 6307;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 109;
        test_state <= test_b1_S6324;
      end
      test_b1_S6324: begin
        IMAGE_addr <= 6308;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 112;
        test_state <= test_b1_S6325;
      end
      test_b1_S6325: begin
        IMAGE_addr <= 6309;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 108;
        test_state <= test_b1_S6326;
      end
      test_b1_S6326: begin
        IMAGE_addr <= 6310;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S6327;
      end
      test_b1_S6327: begin
        IMAGE_addr <= 6311;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6328;
      end
      test_b1_S6328: begin
        IMAGE_addr <= 6312;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S6329;
      end
      test_b1_S6329: begin
        IMAGE_addr <= 6313;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6317;
        test_state <= test_b1_S6330;
      end
      test_b1_S6330: begin
        IMAGE_addr <= 6314;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S6331;
      end
      test_b1_S6331: begin
        IMAGE_addr <= 6315;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 359;
        test_state <= test_b1_S6332;
      end
      test_b1_S6332: begin
        IMAGE_addr <= 6316;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6333;
      end
      test_b1_S6333: begin
        IMAGE_addr <= 6317;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6334;
      end
      test_b1_S6334: begin
        IMAGE_addr <= 6318;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S6335;
      end
      test_b1_S6335: begin
        IMAGE_addr <= 6319;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4066;
        test_state <= test_b1_S6336;
      end
      test_b1_S6336: begin
        IMAGE_addr <= 6320;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6337;
      end
      test_b1_S6337: begin
        IMAGE_addr <= 6321;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6338;
      end
      test_b1_S6338: begin
        IMAGE_addr <= 6322;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S6339;
      end
      test_b1_S6339: begin
        IMAGE_addr <= 6323;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6343;
        test_state <= test_b1_S6340;
      end
      test_b1_S6340: begin
        IMAGE_addr <= 6324;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6341;
      end
      test_b1_S6341: begin
        IMAGE_addr <= 6325;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 344;
        test_state <= test_b1_S6342;
      end
      test_b1_S6342: begin
        IMAGE_addr <= 6326;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 155;
        test_state <= test_b1_S6343;
      end
      test_b1_S6343: begin
        IMAGE_addr <= 6327;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6344;
      end
      test_b1_S6344: begin
        IMAGE_addr <= 6328;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6097;
        test_state <= test_b1_S6345;
      end
      test_b1_S6345: begin
        IMAGE_addr <= 6329;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S6346;
      end
      test_b1_S6346: begin
        IMAGE_addr <= 6330;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S6347;
      end
      test_b1_S6347: begin
        IMAGE_addr <= 6331;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6335;
        test_state <= test_b1_S6348;
      end
      test_b1_S6348: begin
        IMAGE_addr <= 6332;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6271;
        test_state <= test_b1_S6349;
      end
      test_b1_S6349: begin
        IMAGE_addr <= 6333;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S6350;
      end
      test_b1_S6350: begin
        IMAGE_addr <= 6334;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6351;
      end
      test_b1_S6351: begin
        IMAGE_addr <= 6335;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6352;
      end
      test_b1_S6352: begin
        IMAGE_addr <= 6336;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6312;
        test_state <= test_b1_S6353;
      end
      test_b1_S6353: begin
        IMAGE_addr <= 6337;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 732;
        test_state <= test_b1_S6354;
      end
      test_b1_S6354: begin
        IMAGE_addr <= 6338;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6355;
      end
      test_b1_S6355: begin
        IMAGE_addr <= 6339;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 344;
        test_state <= test_b1_S6356;
      end
      test_b1_S6356: begin
        IMAGE_addr <= 6340;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 147;
        test_state <= test_b1_S6357;
      end
      test_b1_S6357: begin
        IMAGE_addr <= 6341;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 345;
        test_state <= test_b1_S6358;
      end
      test_b1_S6358: begin
        IMAGE_addr <= 6342;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6359;
      end
      test_b1_S6359: begin
        IMAGE_addr <= 6343;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6084;
        test_state <= test_b1_S6360;
      end
      test_b1_S6360: begin
        IMAGE_addr <= 6344;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S6361;
      end
      test_b1_S6361: begin
        IMAGE_addr <= 6345;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6352;
        test_state <= test_b1_S6362;
      end
      test_b1_S6362: begin
        IMAGE_addr <= 6346;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 100;
        test_state <= test_b1_S6363;
      end
      test_b1_S6363: begin
        IMAGE_addr <= 6347;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S6364;
      end
      test_b1_S6364: begin
        IMAGE_addr <= 6348;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 112;
        test_state <= test_b1_S6365;
      end
      test_b1_S6365: begin
        IMAGE_addr <= 6349;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S6366;
      end
      test_b1_S6366: begin
        IMAGE_addr <= 6350;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 104;
        test_state <= test_b1_S6367;
      end
      test_b1_S6367: begin
        IMAGE_addr <= 6351;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6368;
      end
      test_b1_S6368: begin
        IMAGE_addr <= 6352;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6369;
      end
      test_b1_S6369: begin
        IMAGE_addr <= 6353;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6370;
      end
      test_b1_S6370: begin
        IMAGE_addr <= 6354;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6371;
      end
      test_b1_S6371: begin
        IMAGE_addr <= 6355;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4294967291;
        test_state <= test_b1_S6372;
      end
      test_b1_S6372: begin
        IMAGE_addr <= 6356;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6373;
      end
      test_b1_S6373: begin
        IMAGE_addr <= 6357;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5;
        test_state <= test_b1_S6374;
      end
      test_b1_S6374: begin
        IMAGE_addr <= 6358;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 29;
        test_state <= test_b1_S6375;
      end
      test_b1_S6375: begin
        IMAGE_addr <= 6359;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 122;
        test_state <= test_b1_S6376;
      end
      test_b1_S6376: begin
        IMAGE_addr <= 6360;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6377;
      end
      test_b1_S6377: begin
        IMAGE_addr <= 6361;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5;
        test_state <= test_b1_S6378;
      end
      test_b1_S6378: begin
        IMAGE_addr <= 6362;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 28;
        test_state <= test_b1_S6379;
      end
      test_b1_S6379: begin
        IMAGE_addr <= 6363;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6380;
      end
      test_b1_S6380: begin
        IMAGE_addr <= 6364;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6381;
      end
      test_b1_S6381: begin
        IMAGE_addr <= 6365;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6343;
        test_state <= test_b1_S6382;
      end
      test_b1_S6382: begin
        IMAGE_addr <= 6366;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S6383;
      end
      test_b1_S6383: begin
        IMAGE_addr <= 6367;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6374;
        test_state <= test_b1_S6384;
      end
      test_b1_S6384: begin
        IMAGE_addr <= 6368;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S6385;
      end
      test_b1_S6385: begin
        IMAGE_addr <= 6369;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S6386;
      end
      test_b1_S6386: begin
        IMAGE_addr <= 6370;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S6387;
      end
      test_b1_S6387: begin
        IMAGE_addr <= 6371;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S6388;
      end
      test_b1_S6388: begin
        IMAGE_addr <= 6372;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S6389;
      end
      test_b1_S6389: begin
        IMAGE_addr <= 6373;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6390;
      end
      test_b1_S6390: begin
        IMAGE_addr <= 6374;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6391;
      end
      test_b1_S6391: begin
        IMAGE_addr <= 6375;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6392;
      end
      test_b1_S6392: begin
        IMAGE_addr <= 6376;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6352;
        test_state <= test_b1_S6393;
      end
      test_b1_S6393: begin
        IMAGE_addr <= 6377;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 25;
        test_state <= test_b1_S6394;
      end
      test_b1_S6394: begin
        IMAGE_addr <= 6378;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 27;
        test_state <= test_b1_S6395;
      end
      test_b1_S6395: begin
        IMAGE_addr <= 6379;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2577;
        test_state <= test_b1_S6396;
      end
      test_b1_S6396: begin
        IMAGE_addr <= 6380;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8;
        test_state <= test_b1_S6397;
      end
      test_b1_S6397: begin
        IMAGE_addr <= 6381;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6377;
        test_state <= test_b1_S6398;
      end
      test_b1_S6398: begin
        IMAGE_addr <= 6382;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6399;
      end
      test_b1_S6399: begin
        IMAGE_addr <= 6383;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6400;
      end
      test_b1_S6400: begin
        IMAGE_addr <= 6384;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6365;
        test_state <= test_b1_S6401;
      end
      test_b1_S6401: begin
        IMAGE_addr <= 6385;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S6402;
      end
      test_b1_S6402: begin
        IMAGE_addr <= 6386;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6392;
        test_state <= test_b1_S6403;
      end
      test_b1_S6403: begin
        IMAGE_addr <= 6387;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 40;
        test_state <= test_b1_S6404;
      end
      test_b1_S6404: begin
        IMAGE_addr <= 6388;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 46;
        test_state <= test_b1_S6405;
      end
      test_b1_S6405: begin
        IMAGE_addr <= 6389;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S6406;
      end
      test_b1_S6406: begin
        IMAGE_addr <= 6390;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 41;
        test_state <= test_b1_S6407;
      end
      test_b1_S6407: begin
        IMAGE_addr <= 6391;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6408;
      end
      test_b1_S6408: begin
        IMAGE_addr <= 6392;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 25;
        test_state <= test_b1_S6409;
      end
      test_b1_S6409: begin
        IMAGE_addr <= 6393;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 27;
        test_state <= test_b1_S6410;
      end
      test_b1_S6410: begin
        IMAGE_addr <= 6394;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S6411;
      end
      test_b1_S6411: begin
        IMAGE_addr <= 6395;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5;
        test_state <= test_b1_S6412;
      end
      test_b1_S6412: begin
        IMAGE_addr <= 6396;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6392;
        test_state <= test_b1_S6413;
      end
      test_b1_S6413: begin
        IMAGE_addr <= 6397;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6;
        test_state <= test_b1_S6414;
      end
      test_b1_S6414: begin
        IMAGE_addr <= 6398;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S6415;
      end
      test_b1_S6415: begin
        IMAGE_addr <= 6399;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4689;
        test_state <= test_b1_S6416;
      end
      test_b1_S6416: begin
        IMAGE_addr <= 6400;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4674;
        test_state <= test_b1_S6417;
      end
      test_b1_S6417: begin
        IMAGE_addr <= 6401;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6418;
      end
      test_b1_S6418: begin
        IMAGE_addr <= 6402;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6419;
      end
      test_b1_S6419: begin
        IMAGE_addr <= 6403;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6365;
        test_state <= test_b1_S6420;
      end
      test_b1_S6420: begin
        IMAGE_addr <= 6404;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S6421;
      end
      test_b1_S6421: begin
        IMAGE_addr <= 6405;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6409;
        test_state <= test_b1_S6422;
      end
      test_b1_S6422: begin
        IMAGE_addr <= 6406;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 46;
        test_state <= test_b1_S6423;
      end
      test_b1_S6423: begin
        IMAGE_addr <= 6407;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S6424;
      end
      test_b1_S6424: begin
        IMAGE_addr <= 6408;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6425;
      end
      test_b1_S6425: begin
        IMAGE_addr <= 6409;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6426;
      end
      test_b1_S6426: begin
        IMAGE_addr <= 6410;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6427;
      end
      test_b1_S6427: begin
        IMAGE_addr <= 6411;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6352;
        test_state <= test_b1_S6428;
      end
      test_b1_S6428: begin
        IMAGE_addr <= 6412;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S6429;
      end
      test_b1_S6429: begin
        IMAGE_addr <= 6413;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6428;
        test_state <= test_b1_S6430;
      end
      test_b1_S6430: begin
        IMAGE_addr <= 6414;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8;
        test_state <= test_b1_S6431;
      end
      test_b1_S6431: begin
        IMAGE_addr <= 6415;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6424;
        test_state <= test_b1_S6432;
      end
      test_b1_S6432: begin
        IMAGE_addr <= 6416;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 92;
        test_state <= test_b1_S6433;
      end
      test_b1_S6433: begin
        IMAGE_addr <= 6417;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 110;
        test_state <= test_b1_S6434;
      end
      test_b1_S6434: begin
        IMAGE_addr <= 6418;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 60;
        test_state <= test_b1_S6435;
      end
      test_b1_S6435: begin
        IMAGE_addr <= 6419;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 37;
        test_state <= test_b1_S6436;
      end
      test_b1_S6436: begin
        IMAGE_addr <= 6420;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 100;
        test_state <= test_b1_S6437;
      end
      test_b1_S6437: begin
        IMAGE_addr <= 6421;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 62;
        test_state <= test_b1_S6438;
      end
      test_b1_S6438: begin
        IMAGE_addr <= 6422;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 32;
        test_state <= test_b1_S6439;
      end
      test_b1_S6439: begin
        IMAGE_addr <= 6423;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6440;
      end
      test_b1_S6440: begin
        IMAGE_addr <= 6424;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6441;
      end
      test_b1_S6441: begin
        IMAGE_addr <= 6425;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6416;
        test_state <= test_b1_S6442;
      end
      test_b1_S6442: begin
        IMAGE_addr <= 6426;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 391;
        test_state <= test_b1_S6443;
      end
      test_b1_S6443: begin
        IMAGE_addr <= 6427;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6444;
      end
      test_b1_S6444: begin
        IMAGE_addr <= 6428;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 774;
        test_state <= test_b1_S6445;
      end
      test_b1_S6445: begin
        IMAGE_addr <= 6429;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6392;
        test_state <= test_b1_S6446;
      end
      test_b1_S6446: begin
        IMAGE_addr <= 6430;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6447;
      end
      test_b1_S6447: begin
        IMAGE_addr <= 6431;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6448;
      end
      test_b1_S6448: begin
        IMAGE_addr <= 6432;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6403;
        test_state <= test_b1_S6449;
      end
      test_b1_S6449: begin
        IMAGE_addr <= 6433;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S6450;
      end
      test_b1_S6450: begin
        IMAGE_addr <= 6434;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6440;
        test_state <= test_b1_S6451;
      end
      test_b1_S6451: begin
        IMAGE_addr <= 6435;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 108;
        test_state <= test_b1_S6452;
      end
      test_b1_S6452: begin
        IMAGE_addr <= 6436;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S6453;
      end
      test_b1_S6453: begin
        IMAGE_addr <= 6437;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S6454;
      end
      test_b1_S6454: begin
        IMAGE_addr <= 6438;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S6455;
      end
      test_b1_S6455: begin
        IMAGE_addr <= 6439;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6456;
      end
      test_b1_S6456: begin
        IMAGE_addr <= 6440;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S6457;
      end
      test_b1_S6457: begin
        IMAGE_addr <= 6441;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6446;
        test_state <= test_b1_S6458;
      end
      test_b1_S6458: begin
        IMAGE_addr <= 6442;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 589;
        test_state <= test_b1_S6459;
      end
      test_b1_S6459: begin
        IMAGE_addr <= 6443;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 391;
        test_state <= test_b1_S6460;
      end
      test_b1_S6460: begin
        IMAGE_addr <= 6444;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4674;
        test_state <= test_b1_S6461;
      end
      test_b1_S6461: begin
        IMAGE_addr <= 6445;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6462;
      end
      test_b1_S6462: begin
        IMAGE_addr <= 6446;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6463;
      end
      test_b1_S6463: begin
        IMAGE_addr <= 6447;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S6464;
      end
      test_b1_S6464: begin
        IMAGE_addr <= 6448;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4066;
        test_state <= test_b1_S6465;
      end
      test_b1_S6465: begin
        IMAGE_addr <= 6449;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6466;
      end
      test_b1_S6466: begin
        IMAGE_addr <= 6450;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6467;
      end
      test_b1_S6467: begin
        IMAGE_addr <= 6451;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6432;
        test_state <= test_b1_S6468;
      end
      test_b1_S6468: begin
        IMAGE_addr <= 6452;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S6469;
      end
      test_b1_S6469: begin
        IMAGE_addr <= 6453;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6461;
        test_state <= test_b1_S6470;
      end
      test_b1_S6470: begin
        IMAGE_addr <= 6454;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 111;
        test_state <= test_b1_S6471;
      end
      test_b1_S6471: begin
        IMAGE_addr <= 6455;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S6472;
      end
      test_b1_S6472: begin
        IMAGE_addr <= 6456;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 104;
        test_state <= test_b1_S6473;
      end
      test_b1_S6473: begin
        IMAGE_addr <= 6457;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S6474;
      end
      test_b1_S6474: begin
        IMAGE_addr <= 6458;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S6475;
      end
      test_b1_S6475: begin
        IMAGE_addr <= 6459;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S6476;
      end
      test_b1_S6476: begin
        IMAGE_addr <= 6460;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6477;
      end
      test_b1_S6477: begin
        IMAGE_addr <= 6461;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6478;
      end
      test_b1_S6478: begin
        IMAGE_addr <= 6462;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4813;
        test_state <= test_b1_S6479;
      end
      test_b1_S6479: begin
        IMAGE_addr <= 6463;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S6480;
      end
      test_b1_S6480: begin
        IMAGE_addr <= 6464;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 25;
        test_state <= test_b1_S6481;
      end
      test_b1_S6481: begin
        IMAGE_addr <= 6465;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 371;
        test_state <= test_b1_S6482;
      end
      test_b1_S6482: begin
        IMAGE_addr <= 6466;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S6483;
      end
      test_b1_S6483: begin
        IMAGE_addr <= 6467;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6484;
      end
      test_b1_S6484: begin
        IMAGE_addr <= 6468;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4813;
        test_state <= test_b1_S6485;
      end
      test_b1_S6485: begin
        IMAGE_addr <= 6469;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 16;
        test_state <= test_b1_S6486;
      end
      test_b1_S6486: begin
        IMAGE_addr <= 6470;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6440;
        test_state <= test_b1_S6487;
      end
      test_b1_S6487: begin
        IMAGE_addr <= 6471;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 27;
        test_state <= test_b1_S6488;
      end
      test_b1_S6488: begin
        IMAGE_addr <= 6472;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8;
        test_state <= test_b1_S6489;
      end
      test_b1_S6489: begin
        IMAGE_addr <= 6473;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6464;
        test_state <= test_b1_S6490;
      end
      test_b1_S6490: begin
        IMAGE_addr <= 6474;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6491;
      end
      test_b1_S6491: begin
        IMAGE_addr <= 6475;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6492;
      end
      test_b1_S6492: begin
        IMAGE_addr <= 6476;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6403;
        test_state <= test_b1_S6493;
      end
      test_b1_S6493: begin
        IMAGE_addr <= 6477;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S6494;
      end
      test_b1_S6494: begin
        IMAGE_addr <= 6478;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6485;
        test_state <= test_b1_S6495;
      end
      test_b1_S6495: begin
        IMAGE_addr <= 6479;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 119;
        test_state <= test_b1_S6496;
      end
      test_b1_S6496: begin
        IMAGE_addr <= 6480;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 111;
        test_state <= test_b1_S6497;
      end
      test_b1_S6497: begin
        IMAGE_addr <= 6481;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S6498;
      end
      test_b1_S6498: begin
        IMAGE_addr <= 6482;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 100;
        test_state <= test_b1_S6499;
      end
      test_b1_S6499: begin
        IMAGE_addr <= 6483;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S6500;
      end
      test_b1_S6500: begin
        IMAGE_addr <= 6484;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6501;
      end
      test_b1_S6501: begin
        IMAGE_addr <= 6485;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6502;
      end
      test_b1_S6502: begin
        IMAGE_addr <= 6486;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6503;
      end
      test_b1_S6503: begin
        IMAGE_addr <= 6487;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 371;
        test_state <= test_b1_S6504;
      end
      test_b1_S6504: begin
        IMAGE_addr <= 6488;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6505;
      end
      test_b1_S6505: begin
        IMAGE_addr <= 6489;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6097;
        test_state <= test_b1_S6506;
      end
      test_b1_S6506: begin
        IMAGE_addr <= 6490;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S6507;
      end
      test_b1_S6507: begin
        IMAGE_addr <= 6491;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S6508;
      end
      test_b1_S6508: begin
        IMAGE_addr <= 6492;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6500;
        test_state <= test_b1_S6509;
      end
      test_b1_S6509: begin
        IMAGE_addr <= 6493;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 155;
        test_state <= test_b1_S6510;
      end
      test_b1_S6510: begin
        IMAGE_addr <= 6494;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6461;
        test_state <= test_b1_S6511;
      end
      test_b1_S6511: begin
        IMAGE_addr <= 6495;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 371;
        test_state <= test_b1_S6512;
      end
      test_b1_S6512: begin
        IMAGE_addr <= 6496;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6513;
      end
      test_b1_S6513: begin
        IMAGE_addr <= 6497;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S6514;
      end
      test_b1_S6514: begin
        IMAGE_addr <= 6498;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6440;
        test_state <= test_b1_S6515;
      end
      test_b1_S6515: begin
        IMAGE_addr <= 6499;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6516;
      end
      test_b1_S6516: begin
        IMAGE_addr <= 6500;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3673;
        test_state <= test_b1_S6517;
      end
      test_b1_S6517: begin
        IMAGE_addr <= 6501;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6518;
      end
      test_b1_S6518: begin
        IMAGE_addr <= 6502;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6519;
      end
      test_b1_S6519: begin
        IMAGE_addr <= 6503;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6476;
        test_state <= test_b1_S6520;
      end
      test_b1_S6520: begin
        IMAGE_addr <= 6504;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S6521;
      end
      test_b1_S6521: begin
        IMAGE_addr <= 6505;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6511;
        test_state <= test_b1_S6522;
      end
      test_b1_S6522: begin
        IMAGE_addr <= 6506;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S6523;
      end
      test_b1_S6523: begin
        IMAGE_addr <= 6507;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S6524;
      end
      test_b1_S6524: begin
        IMAGE_addr <= 6508;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 118;
        test_state <= test_b1_S6525;
      end
      test_b1_S6525: begin
        IMAGE_addr <= 6509;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S6526;
      end
      test_b1_S6526: begin
        IMAGE_addr <= 6510;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6527;
      end
      test_b1_S6527: begin
        IMAGE_addr <= 6511;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6528;
      end
      test_b1_S6528: begin
        IMAGE_addr <= 6512;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6529;
      end
      test_b1_S6529: begin
        IMAGE_addr <= 6513;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6530;
      end
      test_b1_S6530: begin
        IMAGE_addr <= 6514;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6531;
      end
      test_b1_S6531: begin
        IMAGE_addr <= 6515;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6532;
      end
      test_b1_S6532: begin
        IMAGE_addr <= 6516;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S6533;
      end
      test_b1_S6533: begin
        IMAGE_addr <= 6517;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 29;
        test_state <= test_b1_S6534;
      end
      test_b1_S6534: begin
        IMAGE_addr <= 6518;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 122;
        test_state <= test_b1_S6535;
      end
      test_b1_S6535: begin
        IMAGE_addr <= 6519;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6536;
      end
      test_b1_S6536: begin
        IMAGE_addr <= 6520;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6537;
      end
      test_b1_S6537: begin
        IMAGE_addr <= 6521;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6503;
        test_state <= test_b1_S6538;
      end
      test_b1_S6538: begin
        IMAGE_addr <= 6522;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S6539;
      end
      test_b1_S6539: begin
        IMAGE_addr <= 6523;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6528;
        test_state <= test_b1_S6540;
      end
      test_b1_S6540: begin
        IMAGE_addr <= 6524;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 98;
        test_state <= test_b1_S6541;
      end
      test_b1_S6541: begin
        IMAGE_addr <= 6525;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 121;
        test_state <= test_b1_S6542;
      end
      test_b1_S6542: begin
        IMAGE_addr <= 6526;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S6543;
      end
      test_b1_S6543: begin
        IMAGE_addr <= 6527;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6544;
      end
      test_b1_S6544: begin
        IMAGE_addr <= 6528;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6545;
      end
      test_b1_S6545: begin
        IMAGE_addr <= 6529;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6546;
      end
      test_b1_S6546: begin
        IMAGE_addr <= 6530;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 371;
        test_state <= test_b1_S6547;
      end
      test_b1_S6547: begin
        IMAGE_addr <= 6531;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6548;
      end
      test_b1_S6548: begin
        IMAGE_addr <= 6532;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4294967287;
        test_state <= test_b1_S6549;
      end
      test_b1_S6549: begin
        IMAGE_addr <= 6533;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6550;
      end
      test_b1_S6550: begin
        IMAGE_addr <= 6534;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5;
        test_state <= test_b1_S6551;
      end
      test_b1_S6551: begin
        IMAGE_addr <= 6535;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 29;
        test_state <= test_b1_S6552;
      end
      test_b1_S6552: begin
        IMAGE_addr <= 6536;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 122;
        test_state <= test_b1_S6553;
      end
      test_b1_S6553: begin
        IMAGE_addr <= 6537;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6554;
      end
      test_b1_S6554: begin
        IMAGE_addr <= 6538;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6555;
      end
      test_b1_S6555: begin
        IMAGE_addr <= 6539;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6521;
        test_state <= test_b1_S6556;
      end
      test_b1_S6556: begin
        IMAGE_addr <= 6540;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S6557;
      end
      test_b1_S6557: begin
        IMAGE_addr <= 6541;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6551;
        test_state <= test_b1_S6558;
      end
      test_b1_S6558: begin
        IMAGE_addr <= 6542;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 103;
        test_state <= test_b1_S6559;
      end
      test_b1_S6559: begin
        IMAGE_addr <= 6543;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S6560;
      end
      test_b1_S6560: begin
        IMAGE_addr <= 6544;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S6561;
      end
      test_b1_S6561: begin
        IMAGE_addr <= 6545;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 84;
        test_state <= test_b1_S6562;
      end
      test_b1_S6562: begin
        IMAGE_addr <= 6546;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 111;
        test_state <= test_b1_S6563;
      end
      test_b1_S6563: begin
        IMAGE_addr <= 6547;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 107;
        test_state <= test_b1_S6564;
      end
      test_b1_S6564: begin
        IMAGE_addr <= 6548;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S6565;
      end
      test_b1_S6565: begin
        IMAGE_addr <= 6549;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 110;
        test_state <= test_b1_S6566;
      end
      test_b1_S6566: begin
        IMAGE_addr <= 6550;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6567;
      end
      test_b1_S6567: begin
        IMAGE_addr <= 6551;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6568;
      end
      test_b1_S6568: begin
        IMAGE_addr <= 6552;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6569;
      end
      test_b1_S6569: begin
        IMAGE_addr <= 6553;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6570;
      end
      test_b1_S6570: begin
        IMAGE_addr <= 6554;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 32;
        test_state <= test_b1_S6571;
      end
      test_b1_S6571: begin
        IMAGE_addr <= 6555;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 562;
        test_state <= test_b1_S6572;
      end
      test_b1_S6572: begin
        IMAGE_addr <= 6556;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 400;
        test_state <= test_b1_S6573;
      end
      test_b1_S6573: begin
        IMAGE_addr <= 6557;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5792;
        test_state <= test_b1_S6574;
      end
      test_b1_S6574: begin
        IMAGE_addr <= 6558;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6575;
      end
      test_b1_S6575: begin
        IMAGE_addr <= 6559;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6576;
      end
      test_b1_S6576: begin
        IMAGE_addr <= 6560;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6539;
        test_state <= test_b1_S6577;
      end
      test_b1_S6577: begin
        IMAGE_addr <= 6561;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S6578;
      end
      test_b1_S6578: begin
        IMAGE_addr <= 6562;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6573;
        test_state <= test_b1_S6579;
      end
      test_b1_S6579: begin
        IMAGE_addr <= 6563;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 103;
        test_state <= test_b1_S6580;
      end
      test_b1_S6580: begin
        IMAGE_addr <= 6564;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S6581;
      end
      test_b1_S6581: begin
        IMAGE_addr <= 6565;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S6582;
      end
      test_b1_S6582: begin
        IMAGE_addr <= 6566;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 78;
        test_state <= test_b1_S6583;
      end
      test_b1_S6583: begin
        IMAGE_addr <= 6567;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 117;
        test_state <= test_b1_S6584;
      end
      test_b1_S6584: begin
        IMAGE_addr <= 6568;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 109;
        test_state <= test_b1_S6585;
      end
      test_b1_S6585: begin
        IMAGE_addr <= 6569;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 98;
        test_state <= test_b1_S6586;
      end
      test_b1_S6586: begin
        IMAGE_addr <= 6570;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S6587;
      end
      test_b1_S6587: begin
        IMAGE_addr <= 6571;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S6588;
      end
      test_b1_S6588: begin
        IMAGE_addr <= 6572;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6589;
      end
      test_b1_S6589: begin
        IMAGE_addr <= 6573;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6590;
      end
      test_b1_S6590: begin
        IMAGE_addr <= 6574;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6591;
      end
      test_b1_S6591: begin
        IMAGE_addr <= 6575;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6551;
        test_state <= test_b1_S6592;
      end
      test_b1_S6592: begin
        IMAGE_addr <= 6576;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1056;
        test_state <= test_b1_S6593;
      end
      test_b1_S6593: begin
        IMAGE_addr <= 6577;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6594;
      end
      test_b1_S6594: begin
        IMAGE_addr <= 6578;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6595;
      end
      test_b1_S6595: begin
        IMAGE_addr <= 6579;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6560;
        test_state <= test_b1_S6596;
      end
      test_b1_S6596: begin
        IMAGE_addr <= 6580;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S6597;
      end
      test_b1_S6597: begin
        IMAGE_addr <= 6581;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6591;
        test_state <= test_b1_S6598;
      end
      test_b1_S6598: begin
        IMAGE_addr <= 6582;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 58;
        test_state <= test_b1_S6599;
      end
      test_b1_S6599: begin
        IMAGE_addr <= 6583;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S6600;
      end
      test_b1_S6600: begin
        IMAGE_addr <= 6584;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 110;
        test_state <= test_b1_S6601;
      end
      test_b1_S6601: begin
        IMAGE_addr <= 6585;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 99;
        test_state <= test_b1_S6602;
      end
      test_b1_S6602: begin
        IMAGE_addr <= 6586;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 108;
        test_state <= test_b1_S6603;
      end
      test_b1_S6603: begin
        IMAGE_addr <= 6587;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 117;
        test_state <= test_b1_S6604;
      end
      test_b1_S6604: begin
        IMAGE_addr <= 6588;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 100;
        test_state <= test_b1_S6605;
      end
      test_b1_S6605: begin
        IMAGE_addr <= 6589;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S6606;
      end
      test_b1_S6606: begin
        IMAGE_addr <= 6590;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6607;
      end
      test_b1_S6607: begin
        IMAGE_addr <= 6591;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6608;
      end
      test_b1_S6608: begin
        IMAGE_addr <= 6592;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6609;
      end
      test_b1_S6609: begin
        IMAGE_addr <= 6593;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6610;
      end
      test_b1_S6610: begin
        IMAGE_addr <= 6594;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S6611;
      end
      test_b1_S6611: begin
        IMAGE_addr <= 6595;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6612;
      end
      test_b1_S6612: begin
        IMAGE_addr <= 6596;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S6613;
      end
      test_b1_S6613: begin
        IMAGE_addr <= 6597;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 29;
        test_state <= test_b1_S6614;
      end
      test_b1_S6614: begin
        IMAGE_addr <= 6598;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 122;
        test_state <= test_b1_S6615;
      end
      test_b1_S6615: begin
        IMAGE_addr <= 6599;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6616;
      end
      test_b1_S6616: begin
        IMAGE_addr <= 6600;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6617;
      end
      test_b1_S6617: begin
        IMAGE_addr <= 6601;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6579;
        test_state <= test_b1_S6618;
      end
      test_b1_S6618: begin
        IMAGE_addr <= 6602;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S6619;
      end
      test_b1_S6619: begin
        IMAGE_addr <= 6603;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6612;
        test_state <= test_b1_S6620;
      end
      test_b1_S6620: begin
        IMAGE_addr <= 6604;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S6621;
      end
      test_b1_S6621: begin
        IMAGE_addr <= 6605;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 110;
        test_state <= test_b1_S6622;
      end
      test_b1_S6622: begin
        IMAGE_addr <= 6606;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 99;
        test_state <= test_b1_S6623;
      end
      test_b1_S6623: begin
        IMAGE_addr <= 6607;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 108;
        test_state <= test_b1_S6624;
      end
      test_b1_S6624: begin
        IMAGE_addr <= 6608;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 117;
        test_state <= test_b1_S6625;
      end
      test_b1_S6625: begin
        IMAGE_addr <= 6609;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 100;
        test_state <= test_b1_S6626;
      end
      test_b1_S6626: begin
        IMAGE_addr <= 6610;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S6627;
      end
      test_b1_S6627: begin
        IMAGE_addr <= 6611;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6628;
      end
      test_b1_S6628: begin
        IMAGE_addr <= 6612;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6629;
      end
      test_b1_S6629: begin
        IMAGE_addr <= 6613;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6630;
      end
      test_b1_S6630: begin
        IMAGE_addr <= 6614;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6551;
        test_state <= test_b1_S6631;
      end
      test_b1_S6631: begin
        IMAGE_addr <= 6615;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6591;
        test_state <= test_b1_S6632;
      end
      test_b1_S6632: begin
        IMAGE_addr <= 6616;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6633;
      end
      test_b1_S6633: begin
        IMAGE_addr <= 6617;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6634;
      end
      test_b1_S6634: begin
        IMAGE_addr <= 6618;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6601;
        test_state <= test_b1_S6635;
      end
      test_b1_S6635: begin
        IMAGE_addr <= 6619;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S6636;
      end
      test_b1_S6636: begin
        IMAGE_addr <= 6620;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6626;
        test_state <= test_b1_S6637;
      end
      test_b1_S6637: begin
        IMAGE_addr <= 6621;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S6638;
      end
      test_b1_S6638: begin
        IMAGE_addr <= 6622;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S6639;
      end
      test_b1_S6639: begin
        IMAGE_addr <= 6623;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 109;
        test_state <= test_b1_S6640;
      end
      test_b1_S6640: begin
        IMAGE_addr <= 6624;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S6641;
      end
      test_b1_S6641: begin
        IMAGE_addr <= 6625;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6642;
      end
      test_b1_S6642: begin
        IMAGE_addr <= 6626;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6643;
      end
      test_b1_S6643: begin
        IMAGE_addr <= 6627;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6644;
      end
      test_b1_S6644: begin
        IMAGE_addr <= 6628;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6645;
      end
      test_b1_S6645: begin
        IMAGE_addr <= 6629;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4294967288;
        test_state <= test_b1_S6646;
      end
      test_b1_S6646: begin
        IMAGE_addr <= 6630;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6647;
      end
      test_b1_S6647: begin
        IMAGE_addr <= 6631;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5;
        test_state <= test_b1_S6648;
      end
      test_b1_S6648: begin
        IMAGE_addr <= 6632;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 29;
        test_state <= test_b1_S6649;
      end
      test_b1_S6649: begin
        IMAGE_addr <= 6633;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 122;
        test_state <= test_b1_S6650;
      end
      test_b1_S6650: begin
        IMAGE_addr <= 6634;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6651;
      end
      test_b1_S6651: begin
        IMAGE_addr <= 6635;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5;
        test_state <= test_b1_S6652;
      end
      test_b1_S6652: begin
        IMAGE_addr <= 6636;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 28;
        test_state <= test_b1_S6653;
      end
      test_b1_S6653: begin
        IMAGE_addr <= 6637;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6654;
      end
      test_b1_S6654: begin
        IMAGE_addr <= 6638;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6655;
      end
      test_b1_S6655: begin
        IMAGE_addr <= 6639;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6618;
        test_state <= test_b1_S6656;
      end
      test_b1_S6656: begin
        IMAGE_addr <= 6640;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S6657;
      end
      test_b1_S6657: begin
        IMAGE_addr <= 6641;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6648;
        test_state <= test_b1_S6658;
      end
      test_b1_S6658: begin
        IMAGE_addr <= 6642;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 100;
        test_state <= test_b1_S6659;
      end
      test_b1_S6659: begin
        IMAGE_addr <= 6643;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S6660;
      end
      test_b1_S6660: begin
        IMAGE_addr <= 6644;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 108;
        test_state <= test_b1_S6661;
      end
      test_b1_S6661: begin
        IMAGE_addr <= 6645;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S6662;
      end
      test_b1_S6662: begin
        IMAGE_addr <= 6646;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 121;
        test_state <= test_b1_S6663;
      end
      test_b1_S6663: begin
        IMAGE_addr <= 6647;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6664;
      end
      test_b1_S6664: begin
        IMAGE_addr <= 6648;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6665;
      end
      test_b1_S6665: begin
        IMAGE_addr <= 6649;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6666;
      end
      test_b1_S6666: begin
        IMAGE_addr <= 6650;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6626;
        test_state <= test_b1_S6667;
      end
      test_b1_S6667: begin
        IMAGE_addr <= 6651;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 16;
        test_state <= test_b1_S6668;
      end
      test_b1_S6668: begin
        IMAGE_addr <= 6652;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S6669;
      end
      test_b1_S6669: begin
        IMAGE_addr <= 6653;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6658;
        test_state <= test_b1_S6670;
      end
      test_b1_S6670: begin
        IMAGE_addr <= 6654;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S6671;
      end
      test_b1_S6671: begin
        IMAGE_addr <= 6655;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6626;
        test_state <= test_b1_S6672;
      end
      test_b1_S6672: begin
        IMAGE_addr <= 6656;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 830;
        test_state <= test_b1_S6673;
      end
      test_b1_S6673: begin
        IMAGE_addr <= 6657;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6674;
      end
      test_b1_S6674: begin
        IMAGE_addr <= 6658;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3433;
        test_state <= test_b1_S6675;
      end
      test_b1_S6675: begin
        IMAGE_addr <= 6659;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S6676;
      end
      test_b1_S6676: begin
        IMAGE_addr <= 6660;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6677;
      end
      test_b1_S6677: begin
        IMAGE_addr <= 6661;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6678;
      end
      test_b1_S6678: begin
        IMAGE_addr <= 6662;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6639;
        test_state <= test_b1_S6679;
      end
      test_b1_S6679: begin
        IMAGE_addr <= 6663;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S6680;
      end
      test_b1_S6680: begin
        IMAGE_addr <= 6664;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6672;
        test_state <= test_b1_S6681;
      end
      test_b1_S6681: begin
        IMAGE_addr <= 6665;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 103;
        test_state <= test_b1_S6682;
      end
      test_b1_S6682: begin
        IMAGE_addr <= 6666;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S6683;
      end
      test_b1_S6683: begin
        IMAGE_addr <= 6667;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S6684;
      end
      test_b1_S6684: begin
        IMAGE_addr <= 6668;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 69;
        test_state <= test_b1_S6685;
      end
      test_b1_S6685: begin
        IMAGE_addr <= 6669;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 110;
        test_state <= test_b1_S6686;
      end
      test_b1_S6686: begin
        IMAGE_addr <= 6670;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 118;
        test_state <= test_b1_S6687;
      end
      test_b1_S6687: begin
        IMAGE_addr <= 6671;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6688;
      end
      test_b1_S6688: begin
        IMAGE_addr <= 6672;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6689;
      end
      test_b1_S6689: begin
        IMAGE_addr <= 6673;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6690;
      end
      test_b1_S6690: begin
        IMAGE_addr <= 6674;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6691;
      end
      test_b1_S6691: begin
        IMAGE_addr <= 6675;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4294967286;
        test_state <= test_b1_S6692;
      end
      test_b1_S6692: begin
        IMAGE_addr <= 6676;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6693;
      end
      test_b1_S6693: begin
        IMAGE_addr <= 6677;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5;
        test_state <= test_b1_S6694;
      end
      test_b1_S6694: begin
        IMAGE_addr <= 6678;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 29;
        test_state <= test_b1_S6695;
      end
      test_b1_S6695: begin
        IMAGE_addr <= 6679;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 122;
        test_state <= test_b1_S6696;
      end
      test_b1_S6696: begin
        IMAGE_addr <= 6680;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6697;
      end
      test_b1_S6697: begin
        IMAGE_addr <= 6681;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6698;
      end
      test_b1_S6698: begin
        IMAGE_addr <= 6682;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6662;
        test_state <= test_b1_S6699;
      end
      test_b1_S6699: begin
        IMAGE_addr <= 6683;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S6700;
      end
      test_b1_S6700: begin
        IMAGE_addr <= 6684;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6691;
        test_state <= test_b1_S6701;
      end
      test_b1_S6701: begin
        IMAGE_addr <= 6685;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 108;
        test_state <= test_b1_S6702;
      end
      test_b1_S6702: begin
        IMAGE_addr <= 6686;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S6703;
      end
      test_b1_S6703: begin
        IMAGE_addr <= 6687;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S6704;
      end
      test_b1_S6704: begin
        IMAGE_addr <= 6688;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S6705;
      end
      test_b1_S6705: begin
        IMAGE_addr <= 6689;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S6706;
      end
      test_b1_S6706: begin
        IMAGE_addr <= 6690;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6707;
      end
      test_b1_S6707: begin
        IMAGE_addr <= 6691;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6708;
      end
      test_b1_S6708: begin
        IMAGE_addr <= 6692;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6709;
      end
      test_b1_S6709: begin
        IMAGE_addr <= 6693;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6;
        test_state <= test_b1_S6710;
      end
      test_b1_S6710: begin
        IMAGE_addr <= 6694;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6;
        test_state <= test_b1_S6711;
      end
      test_b1_S6711: begin
        IMAGE_addr <= 6695;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S6712;
      end
      test_b1_S6712: begin
        IMAGE_addr <= 6696;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5;
        test_state <= test_b1_S6713;
      end
      test_b1_S6713: begin
        IMAGE_addr <= 6697;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5;
        test_state <= test_b1_S6714;
      end
      test_b1_S6714: begin
        IMAGE_addr <= 6698;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6715;
      end
      test_b1_S6715: begin
        IMAGE_addr <= 6699;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6716;
      end
      test_b1_S6716: begin
        IMAGE_addr <= 6700;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6682;
        test_state <= test_b1_S6717;
      end
      test_b1_S6717: begin
        IMAGE_addr <= 6701;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S6718;
      end
      test_b1_S6718: begin
        IMAGE_addr <= 6702;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6708;
        test_state <= test_b1_S6719;
      end
      test_b1_S6719: begin
        IMAGE_addr <= 6703;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 100;
        test_state <= test_b1_S6720;
      end
      test_b1_S6720: begin
        IMAGE_addr <= 6704;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 111;
        test_state <= test_b1_S6721;
      end
      test_b1_S6721: begin
        IMAGE_addr <= 6705;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 99;
        test_state <= test_b1_S6722;
      end
      test_b1_S6722: begin
        IMAGE_addr <= 6706;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 123;
        test_state <= test_b1_S6723;
      end
      test_b1_S6723: begin
        IMAGE_addr <= 6707;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6724;
      end
      test_b1_S6724: begin
        IMAGE_addr <= 6708;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6725;
      end
      test_b1_S6725: begin
        IMAGE_addr <= 6709;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6726;
      end
      test_b1_S6726: begin
        IMAGE_addr <= 6710;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6551;
        test_state <= test_b1_S6727;
      end
      test_b1_S6727: begin
        IMAGE_addr <= 6711;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8;
        test_state <= test_b1_S6728;
      end
      test_b1_S6728: begin
        IMAGE_addr <= 6712;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6718;
        test_state <= test_b1_S6729;
      end
      test_b1_S6729: begin
        IMAGE_addr <= 6713;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 125;
        test_state <= test_b1_S6730;
      end
      test_b1_S6730: begin
        IMAGE_addr <= 6714;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 100;
        test_state <= test_b1_S6731;
      end
      test_b1_S6731: begin
        IMAGE_addr <= 6715;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 111;
        test_state <= test_b1_S6732;
      end
      test_b1_S6732: begin
        IMAGE_addr <= 6716;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 99;
        test_state <= test_b1_S6733;
      end
      test_b1_S6733: begin
        IMAGE_addr <= 6717;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6734;
      end
      test_b1_S6734: begin
        IMAGE_addr <= 6718;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6735;
      end
      test_b1_S6735: begin
        IMAGE_addr <= 6719;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6713;
        test_state <= test_b1_S6736;
      end
      test_b1_S6736: begin
        IMAGE_addr <= 6720;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 838;
        test_state <= test_b1_S6737;
      end
      test_b1_S6737: begin
        IMAGE_addr <= 6721;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 140;
        test_state <= test_b1_S6738;
      end
      test_b1_S6738: begin
        IMAGE_addr <= 6722;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 25;
        test_state <= test_b1_S6739;
      end
      test_b1_S6739: begin
        IMAGE_addr <= 6723;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S6740;
      end
      test_b1_S6740: begin
        IMAGE_addr <= 6724;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8;
        test_state <= test_b1_S6741;
      end
      test_b1_S6741: begin
        IMAGE_addr <= 6725;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6710;
        test_state <= test_b1_S6742;
      end
      test_b1_S6742: begin
        IMAGE_addr <= 6726;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6743;
      end
      test_b1_S6743: begin
        IMAGE_addr <= 6727;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6744;
      end
      test_b1_S6744: begin
        IMAGE_addr <= 6728;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6700;
        test_state <= test_b1_S6745;
      end
      test_b1_S6745: begin
        IMAGE_addr <= 6729;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S6746;
      end
      test_b1_S6746: begin
        IMAGE_addr <= 6730;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6742;
        test_state <= test_b1_S6747;
      end
      test_b1_S6747: begin
        IMAGE_addr <= 6731;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 118;
        test_state <= test_b1_S6748;
      end
      test_b1_S6748: begin
        IMAGE_addr <= 6732;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S6749;
      end
      test_b1_S6749: begin
        IMAGE_addr <= 6733;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S6750;
      end
      test_b1_S6750: begin
        IMAGE_addr <= 6734;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S6751;
      end
      test_b1_S6751: begin
        IMAGE_addr <= 6735;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S6752;
      end
      test_b1_S6752: begin
        IMAGE_addr <= 6736;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 98;
        test_state <= test_b1_S6753;
      end
      test_b1_S6753: begin
        IMAGE_addr <= 6737;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 108;
        test_state <= test_b1_S6754;
      end
      test_b1_S6754: begin
        IMAGE_addr <= 6738;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S6755;
      end
      test_b1_S6755: begin
        IMAGE_addr <= 6739;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S6756;
      end
      test_b1_S6756: begin
        IMAGE_addr <= 6740;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 124;
        test_state <= test_b1_S6757;
      end
      test_b1_S6757: begin
        IMAGE_addr <= 6741;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6758;
      end
      test_b1_S6758: begin
        IMAGE_addr <= 6742;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6759;
      end
      test_b1_S6759: begin
        IMAGE_addr <= 6743;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6760;
      end
      test_b1_S6760: begin
        IMAGE_addr <= 6744;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6551;
        test_state <= test_b1_S6761;
      end
      test_b1_S6761: begin
        IMAGE_addr <= 6745;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8;
        test_state <= test_b1_S6762;
      end
      test_b1_S6762: begin
        IMAGE_addr <= 6746;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6749;
        test_state <= test_b1_S6763;
      end
      test_b1_S6763: begin
        IMAGE_addr <= 6747;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 124;
        test_state <= test_b1_S6764;
      end
      test_b1_S6764: begin
        IMAGE_addr <= 6748;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6765;
      end
      test_b1_S6765: begin
        IMAGE_addr <= 6749;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6766;
      end
      test_b1_S6766: begin
        IMAGE_addr <= 6750;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6747;
        test_state <= test_b1_S6767;
      end
      test_b1_S6767: begin
        IMAGE_addr <= 6751;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 838;
        test_state <= test_b1_S6768;
      end
      test_b1_S6768: begin
        IMAGE_addr <= 6752;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 140;
        test_state <= test_b1_S6769;
      end
      test_b1_S6769: begin
        IMAGE_addr <= 6753;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 25;
        test_state <= test_b1_S6770;
      end
      test_b1_S6770: begin
        IMAGE_addr <= 6754;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S6771;
      end
      test_b1_S6771: begin
        IMAGE_addr <= 6755;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 400;
        test_state <= test_b1_S6772;
      end
      test_b1_S6772: begin
        IMAGE_addr <= 6756;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 596;
        test_state <= test_b1_S6773;
      end
      test_b1_S6773: begin
        IMAGE_addr <= 6757;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6774;
      end
      test_b1_S6774: begin
        IMAGE_addr <= 6758;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6775;
      end
      test_b1_S6775: begin
        IMAGE_addr <= 6759;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 213;
        test_state <= test_b1_S6776;
      end
      test_b1_S6776: begin
        IMAGE_addr <= 6760;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8;
        test_state <= test_b1_S6777;
      end
      test_b1_S6777: begin
        IMAGE_addr <= 6761;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6744;
        test_state <= test_b1_S6778;
      end
      test_b1_S6778: begin
        IMAGE_addr <= 6762;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6779;
      end
      test_b1_S6779: begin
        IMAGE_addr <= 6763;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6780;
      end
      test_b1_S6780: begin
        IMAGE_addr <= 6764;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6728;
        test_state <= test_b1_S6781;
      end
      test_b1_S6781: begin
        IMAGE_addr <= 6765;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S6782;
      end
      test_b1_S6782: begin
        IMAGE_addr <= 6766;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6771;
        test_state <= test_b1_S6783;
      end
      test_b1_S6783: begin
        IMAGE_addr <= 6767;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 112;
        test_state <= test_b1_S6784;
      end
      test_b1_S6784: begin
        IMAGE_addr <= 6768;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 111;
        test_state <= test_b1_S6785;
      end
      test_b1_S6785: begin
        IMAGE_addr <= 6769;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 119;
        test_state <= test_b1_S6786;
      end
      test_b1_S6786: begin
        IMAGE_addr <= 6770;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6787;
      end
      test_b1_S6787: begin
        IMAGE_addr <= 6771;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6788;
      end
      test_b1_S6788: begin
        IMAGE_addr <= 6772;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6789;
      end
      test_b1_S6789: begin
        IMAGE_addr <= 6773;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6790;
      end
      test_b1_S6790: begin
        IMAGE_addr <= 6774;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6791;
      end
      test_b1_S6791: begin
        IMAGE_addr <= 6775;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S6792;
      end
      test_b1_S6792: begin
        IMAGE_addr <= 6776;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S6793;
      end
      test_b1_S6793: begin
        IMAGE_addr <= 6777;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6781;
        test_state <= test_b1_S6794;
      end
      test_b1_S6794: begin
        IMAGE_addr <= 6778;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 132;
        test_state <= test_b1_S6795;
      end
      test_b1_S6795: begin
        IMAGE_addr <= 6779;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 18;
        test_state <= test_b1_S6796;
      end
      test_b1_S6796: begin
        IMAGE_addr <= 6780;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6797;
      end
      test_b1_S6797: begin
        IMAGE_addr <= 6781;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3841;
        test_state <= test_b1_S6798;
      end
      test_b1_S6798: begin
        IMAGE_addr <= 6782;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2577;
        test_state <= test_b1_S6799;
      end
      test_b1_S6799: begin
        IMAGE_addr <= 6783;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6800;
      end
      test_b1_S6800: begin
        IMAGE_addr <= 6784;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6801;
      end
      test_b1_S6801: begin
        IMAGE_addr <= 6785;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6764;
        test_state <= test_b1_S6802;
      end
      test_b1_S6802: begin
        IMAGE_addr <= 6786;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S6803;
      end
      test_b1_S6803: begin
        IMAGE_addr <= 6787;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6792;
        test_state <= test_b1_S6804;
      end
      test_b1_S6804: begin
        IMAGE_addr <= 6788;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S6805;
      end
      test_b1_S6805: begin
        IMAGE_addr <= 6789;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 98;
        test_state <= test_b1_S6806;
      end
      test_b1_S6806: begin
        IMAGE_addr <= 6790;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S6807;
      end
      test_b1_S6807: begin
        IMAGE_addr <= 6791;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6808;
      end
      test_b1_S6808: begin
        IMAGE_addr <= 6792;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6809;
      end
      test_b1_S6809: begin
        IMAGE_addr <= 6793;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6810;
      end
      test_b1_S6810: begin
        IMAGE_addr <= 6794;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S6811;
      end
      test_b1_S6811: begin
        IMAGE_addr <= 6795;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6812;
      end
      test_b1_S6812: begin
        IMAGE_addr <= 6796;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6813;
      end
      test_b1_S6813: begin
        IMAGE_addr <= 6797;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 822;
        test_state <= test_b1_S6814;
      end
      test_b1_S6814: begin
        IMAGE_addr <= 6798;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6815;
      end
      test_b1_S6815: begin
        IMAGE_addr <= 6799;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 176;
        test_state <= test_b1_S6816;
      end
      test_b1_S6816: begin
        IMAGE_addr <= 6800;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 751;
        test_state <= test_b1_S6817;
      end
      test_b1_S6817: begin
        IMAGE_addr <= 6801;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6818;
      end
      test_b1_S6818: begin
        IMAGE_addr <= 6802;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6819;
      end
      test_b1_S6819: begin
        IMAGE_addr <= 6803;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6785;
        test_state <= test_b1_S6820;
      end
      test_b1_S6820: begin
        IMAGE_addr <= 6804;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S6821;
      end
      test_b1_S6821: begin
        IMAGE_addr <= 6805;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6810;
        test_state <= test_b1_S6822;
      end
      test_b1_S6822: begin
        IMAGE_addr <= 6806;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 109;
        test_state <= test_b1_S6823;
      end
      test_b1_S6823: begin
        IMAGE_addr <= 6807;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S6824;
      end
      test_b1_S6824: begin
        IMAGE_addr <= 6808;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 110;
        test_state <= test_b1_S6825;
      end
      test_b1_S6825: begin
        IMAGE_addr <= 6809;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6826;
      end
      test_b1_S6826: begin
        IMAGE_addr <= 6810;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6827;
      end
      test_b1_S6827: begin
        IMAGE_addr <= 6811;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6828;
      end
      test_b1_S6828: begin
        IMAGE_addr <= 6812;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 132;
        test_state <= test_b1_S6829;
      end
      test_b1_S6829: begin
        IMAGE_addr <= 6813;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 132;
        test_state <= test_b1_S6830;
      end
      test_b1_S6830: begin
        IMAGE_addr <= 6814;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 822;
        test_state <= test_b1_S6831;
      end
      test_b1_S6831: begin
        IMAGE_addr <= 6815;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6832;
      end
      test_b1_S6832: begin
        IMAGE_addr <= 6816;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 52;
        test_state <= test_b1_S6833;
      end
      test_b1_S6833: begin
        IMAGE_addr <= 6817;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6834;
      end
      test_b1_S6834: begin
        IMAGE_addr <= 6818;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2577;
        test_state <= test_b1_S6835;
      end
      test_b1_S6835: begin
        IMAGE_addr <= 6819;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 732;
        test_state <= test_b1_S6836;
      end
      test_b1_S6836: begin
        IMAGE_addr <= 6820;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6837;
      end
      test_b1_S6837: begin
        IMAGE_addr <= 6821;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6838;
      end
      test_b1_S6838: begin
        IMAGE_addr <= 6822;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6803;
        test_state <= test_b1_S6839;
      end
      test_b1_S6839: begin
        IMAGE_addr <= 6823;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S6840;
      end
      test_b1_S6840: begin
        IMAGE_addr <= 6824;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6829;
        test_state <= test_b1_S6841;
      end
      test_b1_S6841: begin
        IMAGE_addr <= 6825;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 109;
        test_state <= test_b1_S6842;
      end
      test_b1_S6842: begin
        IMAGE_addr <= 6826;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S6843;
      end
      test_b1_S6843: begin
        IMAGE_addr <= 6827;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 120;
        test_state <= test_b1_S6844;
      end
      test_b1_S6844: begin
        IMAGE_addr <= 6828;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6845;
      end
      test_b1_S6845: begin
        IMAGE_addr <= 6829;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6846;
      end
      test_b1_S6846: begin
        IMAGE_addr <= 6830;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6847;
      end
      test_b1_S6847: begin
        IMAGE_addr <= 6831;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 132;
        test_state <= test_b1_S6848;
      end
      test_b1_S6848: begin
        IMAGE_addr <= 6832;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 132;
        test_state <= test_b1_S6849;
      end
      test_b1_S6849: begin
        IMAGE_addr <= 6833;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 822;
        test_state <= test_b1_S6850;
      end
      test_b1_S6850: begin
        IMAGE_addr <= 6834;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6851;
      end
      test_b1_S6851: begin
        IMAGE_addr <= 6835;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2577;
        test_state <= test_b1_S6852;
      end
      test_b1_S6852: begin
        IMAGE_addr <= 6836;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6853;
      end
      test_b1_S6853: begin
        IMAGE_addr <= 6837;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 52;
        test_state <= test_b1_S6854;
      end
      test_b1_S6854: begin
        IMAGE_addr <= 6838;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 732;
        test_state <= test_b1_S6855;
      end
      test_b1_S6855: begin
        IMAGE_addr <= 6839;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6856;
      end
      test_b1_S6856: begin
        IMAGE_addr <= 6840;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6857;
      end
      test_b1_S6857: begin
        IMAGE_addr <= 6841;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6822;
        test_state <= test_b1_S6858;
      end
      test_b1_S6858: begin
        IMAGE_addr <= 6842;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 310;
        test_state <= test_b1_S6859;
      end
      test_b1_S6859: begin
        IMAGE_addr <= 6843;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6846;
        test_state <= test_b1_S6860;
      end
      test_b1_S6860: begin
        IMAGE_addr <= 6844;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 119;
        test_state <= test_b1_S6861;
      end
      test_b1_S6861: begin
        IMAGE_addr <= 6845;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6862;
      end
      test_b1_S6862: begin
        IMAGE_addr <= 6846;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6863;
      end
      test_b1_S6863: begin
        IMAGE_addr <= 6847;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6841;
        test_state <= test_b1_S6864;
      end
      test_b1_S6864: begin
        IMAGE_addr <= 6848;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 310;
        test_state <= test_b1_S6865;
      end
      test_b1_S6865: begin
        IMAGE_addr <= 6849;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6852;
        test_state <= test_b1_S6866;
      end
      test_b1_S6866: begin
        IMAGE_addr <= 6850;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 122;
        test_state <= test_b1_S6867;
      end
      test_b1_S6867: begin
        IMAGE_addr <= 6851;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6868;
      end
      test_b1_S6868: begin
        IMAGE_addr <= 6852;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6869;
      end
      test_b1_S6869: begin
        IMAGE_addr <= 6853;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6847;
        test_state <= test_b1_S6870;
      end
      test_b1_S6870: begin
        IMAGE_addr <= 6854;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S6871;
      end
      test_b1_S6871: begin
        IMAGE_addr <= 6855;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6863;
        test_state <= test_b1_S6872;
      end
      test_b1_S6872: begin
        IMAGE_addr <= 6856;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S6873;
      end
      test_b1_S6873: begin
        IMAGE_addr <= 6857;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S6874;
      end
      test_b1_S6874: begin
        IMAGE_addr <= 6858;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S6875;
      end
      test_b1_S6875: begin
        IMAGE_addr <= 6859;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 100;
        test_state <= test_b1_S6876;
      end
      test_b1_S6876: begin
        IMAGE_addr <= 6860;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S6877;
      end
      test_b1_S6877: begin
        IMAGE_addr <= 6861;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 63;
        test_state <= test_b1_S6878;
      end
      test_b1_S6878: begin
        IMAGE_addr <= 6862;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6879;
      end
      test_b1_S6879: begin
        IMAGE_addr <= 6863;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6880;
      end
      test_b1_S6880: begin
        IMAGE_addr <= 6864;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6846;
        test_state <= test_b1_S6881;
      end
      test_b1_S6881: begin
        IMAGE_addr <= 6865;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S6882;
      end
      test_b1_S6882: begin
        IMAGE_addr <= 6866;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6883;
      end
      test_b1_S6883: begin
        IMAGE_addr <= 6867;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6852;
        test_state <= test_b1_S6884;
      end
      test_b1_S6884: begin
        IMAGE_addr <= 6868;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S6885;
      end
      test_b1_S6885: begin
        IMAGE_addr <= 6869;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 20;
        test_state <= test_b1_S6886;
      end
      test_b1_S6886: begin
        IMAGE_addr <= 6870;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6887;
      end
      test_b1_S6887: begin
        IMAGE_addr <= 6871;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6888;
      end
      test_b1_S6888: begin
        IMAGE_addr <= 6872;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6853;
        test_state <= test_b1_S6889;
      end
      test_b1_S6889: begin
        IMAGE_addr <= 6873;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S6890;
      end
      test_b1_S6890: begin
        IMAGE_addr <= 6874;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6880;
        test_state <= test_b1_S6891;
      end
      test_b1_S6891: begin
        IMAGE_addr <= 6875;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S6892;
      end
      test_b1_S6892: begin
        IMAGE_addr <= 6876;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S6893;
      end
      test_b1_S6893: begin
        IMAGE_addr <= 6877;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S6894;
      end
      test_b1_S6894: begin
        IMAGE_addr <= 6878;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 100;
        test_state <= test_b1_S6895;
      end
      test_b1_S6895: begin
        IMAGE_addr <= 6879;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6896;
      end
      test_b1_S6896: begin
        IMAGE_addr <= 6880;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6626;
        test_state <= test_b1_S6897;
      end
      test_b1_S6897: begin
        IMAGE_addr <= 6881;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S6898;
      end
      test_b1_S6898: begin
        IMAGE_addr <= 6882;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6890;
        test_state <= test_b1_S6899;
      end
      test_b1_S6899: begin
        IMAGE_addr <= 6883;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6900;
      end
      test_b1_S6900: begin
        IMAGE_addr <= 6884;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 62903;
        test_state <= test_b1_S6901;
      end
      test_b1_S6901: begin
        IMAGE_addr <= 6885;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 20;
        test_state <= test_b1_S6902;
      end
      test_b1_S6902: begin
        IMAGE_addr <= 6886;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6903;
      end
      test_b1_S6903: begin
        IMAGE_addr <= 6887;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6846;
        test_state <= test_b1_S6904;
      end
      test_b1_S6904: begin
        IMAGE_addr <= 6888;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S6905;
      end
      test_b1_S6905: begin
        IMAGE_addr <= 6889;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6906;
      end
      test_b1_S6906: begin
        IMAGE_addr <= 6890;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S6907;
      end
      test_b1_S6907: begin
        IMAGE_addr <= 6891;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6899;
        test_state <= test_b1_S6908;
      end
      test_b1_S6908: begin
        IMAGE_addr <= 6892;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6909;
      end
      test_b1_S6909: begin
        IMAGE_addr <= 6893;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 78578;
        test_state <= test_b1_S6910;
      end
      test_b1_S6910: begin
        IMAGE_addr <= 6894;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 20;
        test_state <= test_b1_S6911;
      end
      test_b1_S6911: begin
        IMAGE_addr <= 6895;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6912;
      end
      test_b1_S6912: begin
        IMAGE_addr <= 6896;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6852;
        test_state <= test_b1_S6913;
      end
      test_b1_S6913: begin
        IMAGE_addr <= 6897;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S6914;
      end
      test_b1_S6914: begin
        IMAGE_addr <= 6898;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6915;
      end
      test_b1_S6915: begin
        IMAGE_addr <= 6899;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3539;
        test_state <= test_b1_S6916;
      end
      test_b1_S6916: begin
        IMAGE_addr <= 6900;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6917;
      end
      test_b1_S6917: begin
        IMAGE_addr <= 6901;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6918;
      end
      test_b1_S6918: begin
        IMAGE_addr <= 6902;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6872;
        test_state <= test_b1_S6919;
      end
      test_b1_S6919: begin
        IMAGE_addr <= 6903;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S6920;
      end
      test_b1_S6920: begin
        IMAGE_addr <= 6904;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6911;
        test_state <= test_b1_S6921;
      end
      test_b1_S6921: begin
        IMAGE_addr <= 6905;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 63;
        test_state <= test_b1_S6922;
      end
      test_b1_S6922: begin
        IMAGE_addr <= 6906;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S6923;
      end
      test_b1_S6923: begin
        IMAGE_addr <= 6907;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S6924;
      end
      test_b1_S6924: begin
        IMAGE_addr <= 6908;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S6925;
      end
      test_b1_S6925: begin
        IMAGE_addr <= 6909;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 100;
        test_state <= test_b1_S6926;
      end
      test_b1_S6926: begin
        IMAGE_addr <= 6910;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6927;
      end
      test_b1_S6927: begin
        IMAGE_addr <= 6911;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6863;
        test_state <= test_b1_S6928;
      end
      test_b1_S6928: begin
        IMAGE_addr <= 6912;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6929;
      end
      test_b1_S6929: begin
        IMAGE_addr <= 6913;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6930;
      end
      test_b1_S6930: begin
        IMAGE_addr <= 6914;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 798;
        test_state <= test_b1_S6931;
      end
      test_b1_S6931: begin
        IMAGE_addr <= 6915;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 140;
        test_state <= test_b1_S6932;
      end
      test_b1_S6932: begin
        IMAGE_addr <= 6916;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 25;
        test_state <= test_b1_S6933;
      end
      test_b1_S6933: begin
        IMAGE_addr <= 6917;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S6934;
      end
      test_b1_S6934: begin
        IMAGE_addr <= 6918;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6880;
        test_state <= test_b1_S6935;
      end
      test_b1_S6935: begin
        IMAGE_addr <= 6919;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8;
        test_state <= test_b1_S6936;
      end
      test_b1_S6936: begin
        IMAGE_addr <= 6920;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6911;
        test_state <= test_b1_S6937;
      end
      test_b1_S6937: begin
        IMAGE_addr <= 6921;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6938;
      end
      test_b1_S6938: begin
        IMAGE_addr <= 6922;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S6939;
      end
      test_b1_S6939: begin
        IMAGE_addr <= 6923;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6902;
        test_state <= test_b1_S6940;
      end
      test_b1_S6940: begin
        IMAGE_addr <= 6924;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S6941;
      end
      test_b1_S6941: begin
        IMAGE_addr <= 6925;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6935;
        test_state <= test_b1_S6942;
      end
      test_b1_S6942: begin
        IMAGE_addr <= 6926;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 40;
        test_state <= test_b1_S6943;
      end
      test_b1_S6943: begin
        IMAGE_addr <= 6927;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S6944;
      end
      test_b1_S6944: begin
        IMAGE_addr <= 6928;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S6945;
      end
      test_b1_S6945: begin
        IMAGE_addr <= 6929;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 110;
        test_state <= test_b1_S6946;
      end
      test_b1_S6946: begin
        IMAGE_addr <= 6930;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 100;
        test_state <= test_b1_S6947;
      end
      test_b1_S6947: begin
        IMAGE_addr <= 6931;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 111;
        test_state <= test_b1_S6948;
      end
      test_b1_S6948: begin
        IMAGE_addr <= 6932;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 109;
        test_state <= test_b1_S6949;
      end
      test_b1_S6949: begin
        IMAGE_addr <= 6933;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 41;
        test_state <= test_b1_S6950;
      end
      test_b1_S6950: begin
        IMAGE_addr <= 6934;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S6951;
      end
      test_b1_S6951: begin
        IMAGE_addr <= 6935;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6952;
      end
      test_b1_S6952: begin
        IMAGE_addr <= 6936;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 36969;
        test_state <= test_b1_S6953;
      end
      test_b1_S6953: begin
        IMAGE_addr <= 6937;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6954;
      end
      test_b1_S6954: begin
        IMAGE_addr <= 6938;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6852;
        test_state <= test_b1_S6955;
      end
      test_b1_S6955: begin
        IMAGE_addr <= 6939;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S6956;
      end
      test_b1_S6956: begin
        IMAGE_addr <= 6940;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6957;
      end
      test_b1_S6957: begin
        IMAGE_addr <= 6941;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 65535;
        test_state <= test_b1_S6958;
      end
      test_b1_S6958: begin
        IMAGE_addr <= 6942;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 20;
        test_state <= test_b1_S6959;
      end
      test_b1_S6959: begin
        IMAGE_addr <= 6943;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 18;
        test_state <= test_b1_S6960;
      end
      test_b1_S6960: begin
        IMAGE_addr <= 6944;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6961;
      end
      test_b1_S6961: begin
        IMAGE_addr <= 6945;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6852;
        test_state <= test_b1_S6962;
      end
      test_b1_S6962: begin
        IMAGE_addr <= 6946;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S6963;
      end
      test_b1_S6963: begin
        IMAGE_addr <= 6947;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6964;
      end
      test_b1_S6964: begin
        IMAGE_addr <= 6948;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 16;
        test_state <= test_b1_S6965;
      end
      test_b1_S6965: begin
        IMAGE_addr <= 6949;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 24;
        test_state <= test_b1_S6966;
      end
      test_b1_S6966: begin
        IMAGE_addr <= 6950;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 16;
        test_state <= test_b1_S6967;
      end
      test_b1_S6967: begin
        IMAGE_addr <= 6951;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6968;
      end
      test_b1_S6968: begin
        IMAGE_addr <= 6952;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6852;
        test_state <= test_b1_S6969;
      end
      test_b1_S6969: begin
        IMAGE_addr <= 6953;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S6970;
      end
      test_b1_S6970: begin
        IMAGE_addr <= 6954;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6971;
      end
      test_b1_S6971: begin
        IMAGE_addr <= 6955;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 18000;
        test_state <= test_b1_S6972;
      end
      test_b1_S6972: begin
        IMAGE_addr <= 6956;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6973;
      end
      test_b1_S6973: begin
        IMAGE_addr <= 6957;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6846;
        test_state <= test_b1_S6974;
      end
      test_b1_S6974: begin
        IMAGE_addr <= 6958;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S6975;
      end
      test_b1_S6975: begin
        IMAGE_addr <= 6959;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6976;
      end
      test_b1_S6976: begin
        IMAGE_addr <= 6960;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 65535;
        test_state <= test_b1_S6977;
      end
      test_b1_S6977: begin
        IMAGE_addr <= 6961;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 20;
        test_state <= test_b1_S6978;
      end
      test_b1_S6978: begin
        IMAGE_addr <= 6962;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 18;
        test_state <= test_b1_S6979;
      end
      test_b1_S6979: begin
        IMAGE_addr <= 6963;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6980;
      end
      test_b1_S6980: begin
        IMAGE_addr <= 6964;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6846;
        test_state <= test_b1_S6981;
      end
      test_b1_S6981: begin
        IMAGE_addr <= 6965;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S6982;
      end
      test_b1_S6982: begin
        IMAGE_addr <= 6966;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6983;
      end
      test_b1_S6983: begin
        IMAGE_addr <= 6967;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 16;
        test_state <= test_b1_S6984;
      end
      test_b1_S6984: begin
        IMAGE_addr <= 6968;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 24;
        test_state <= test_b1_S6985;
      end
      test_b1_S6985: begin
        IMAGE_addr <= 6969;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 16;
        test_state <= test_b1_S6986;
      end
      test_b1_S6986: begin
        IMAGE_addr <= 6970;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6987;
      end
      test_b1_S6987: begin
        IMAGE_addr <= 6971;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6846;
        test_state <= test_b1_S6988;
      end
      test_b1_S6988: begin
        IMAGE_addr <= 6972;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S6989;
      end
      test_b1_S6989: begin
        IMAGE_addr <= 6973;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6990;
      end
      test_b1_S6990: begin
        IMAGE_addr <= 6974;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6852;
        test_state <= test_b1_S6991;
      end
      test_b1_S6991: begin
        IMAGE_addr <= 6975;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S6992;
      end
      test_b1_S6992: begin
        IMAGE_addr <= 6976;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6993;
      end
      test_b1_S6993: begin
        IMAGE_addr <= 6977;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 16;
        test_state <= test_b1_S6994;
      end
      test_b1_S6994: begin
        IMAGE_addr <= 6978;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 23;
        test_state <= test_b1_S6995;
      end
      test_b1_S6995: begin
        IMAGE_addr <= 6979;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S6996;
      end
      test_b1_S6996: begin
        IMAGE_addr <= 6980;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6846;
        test_state <= test_b1_S6997;
      end
      test_b1_S6997: begin
        IMAGE_addr <= 6981;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S6998;
      end
      test_b1_S6998: begin
        IMAGE_addr <= 6982;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 16;
        test_state <= test_b1_S6999;
      end
      test_b1_S6999: begin
        IMAGE_addr <= 6983;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7000;
      end
      test_b1_S7000: begin
        IMAGE_addr <= 6984;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7001;
      end
      test_b1_S7001: begin
        IMAGE_addr <= 6985;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6822;
        test_state <= test_b1_S7002;
      end
      test_b1_S7002: begin
        IMAGE_addr <= 6986;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S7003;
      end
      test_b1_S7003: begin
        IMAGE_addr <= 6987;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6995;
        test_state <= test_b1_S7004;
      end
      test_b1_S7004: begin
        IMAGE_addr <= 6988;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S7005;
      end
      test_b1_S7005: begin
        IMAGE_addr <= 6989;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S7006;
      end
      test_b1_S7006: begin
        IMAGE_addr <= 6990;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 110;
        test_state <= test_b1_S7007;
      end
      test_b1_S7007: begin
        IMAGE_addr <= 6991;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 100;
        test_state <= test_b1_S7008;
      end
      test_b1_S7008: begin
        IMAGE_addr <= 6992;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 111;
        test_state <= test_b1_S7009;
      end
      test_b1_S7009: begin
        IMAGE_addr <= 6993;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 109;
        test_state <= test_b1_S7010;
      end
      test_b1_S7010: begin
        IMAGE_addr <= 6994;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7011;
      end
      test_b1_S7011: begin
        IMAGE_addr <= 6995;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7012;
      end
      test_b1_S7012: begin
        IMAGE_addr <= 6996;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7013;
      end
      test_b1_S7013: begin
        IMAGE_addr <= 6997;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6911;
        test_state <= test_b1_S7014;
      end
      test_b1_S7014: begin
        IMAGE_addr <= 6998;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6935;
        test_state <= test_b1_S7015;
      end
      test_b1_S7015: begin
        IMAGE_addr <= 6999;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6792;
        test_state <= test_b1_S7016;
      end
      test_b1_S7016: begin
        IMAGE_addr <= 7000;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7017;
      end
      test_b1_S7017: begin
        IMAGE_addr <= 7001;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7018;
      end
      test_b1_S7018: begin
        IMAGE_addr <= 7002;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6985;
        test_state <= test_b1_S7019;
      end
      test_b1_S7019: begin
        IMAGE_addr <= 7003;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5034;
        test_state <= test_b1_S7020;
      end
      test_b1_S7020: begin
        IMAGE_addr <= 7004;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7157;
        test_state <= test_b1_S7021;
      end
      test_b1_S7021: begin
        IMAGE_addr <= 7005;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 98;
        test_state <= test_b1_S7022;
      end
      test_b1_S7022: begin
        IMAGE_addr <= 7006;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 117;
        test_state <= test_b1_S7023;
      end
      test_b1_S7023: begin
        IMAGE_addr <= 7007;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 102;
        test_state <= test_b1_S7024;
      end
      test_b1_S7024: begin
        IMAGE_addr <= 7008;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 102;
        test_state <= test_b1_S7025;
      end
      test_b1_S7025: begin
        IMAGE_addr <= 7009;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S7026;
      end
      test_b1_S7026: begin
        IMAGE_addr <= 7010;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S7027;
      end
      test_b1_S7027: begin
        IMAGE_addr <= 7011;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 39;
        test_state <= test_b1_S7028;
      end
      test_b1_S7028: begin
        IMAGE_addr <= 7012;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7029;
      end
      test_b1_S7029: begin
        IMAGE_addr <= 7013;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7030;
      end
      test_b1_S7030: begin
        IMAGE_addr <= 7014;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7031;
      end
      test_b1_S7031: begin
        IMAGE_addr <= 7015;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 306;
        test_state <= test_b1_S7032;
      end
      test_b1_S7032: begin
        IMAGE_addr <= 7016;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4956;
        test_state <= test_b1_S7033;
      end
      test_b1_S7033: begin
        IMAGE_addr <= 7017;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 37;
        test_state <= test_b1_S7034;
      end
      test_b1_S7034: begin
        IMAGE_addr <= 7018;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 37;
        test_state <= test_b1_S7035;
      end
      test_b1_S7035: begin
        IMAGE_addr <= 7019;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7036;
      end
      test_b1_S7036: begin
        IMAGE_addr <= 7020;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7014;
        test_state <= test_b1_S7037;
      end
      test_b1_S7037: begin
        IMAGE_addr <= 7021;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 310;
        test_state <= test_b1_S7038;
      end
      test_b1_S7038: begin
        IMAGE_addr <= 7022;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7030;
        test_state <= test_b1_S7039;
      end
      test_b1_S7039: begin
        IMAGE_addr <= 7023;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 98;
        test_state <= test_b1_S7040;
      end
      test_b1_S7040: begin
        IMAGE_addr <= 7024;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 117;
        test_state <= test_b1_S7041;
      end
      test_b1_S7041: begin
        IMAGE_addr <= 7025;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 102;
        test_state <= test_b1_S7042;
      end
      test_b1_S7042: begin
        IMAGE_addr <= 7026;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 102;
        test_state <= test_b1_S7043;
      end
      test_b1_S7043: begin
        IMAGE_addr <= 7027;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S7044;
      end
      test_b1_S7044: begin
        IMAGE_addr <= 7028;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S7045;
      end
      test_b1_S7045: begin
        IMAGE_addr <= 7029;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7046;
      end
      test_b1_S7046: begin
        IMAGE_addr <= 7030;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7047;
      end
      test_b1_S7047: begin
        IMAGE_addr <= 7031;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7020;
        test_state <= test_b1_S7048;
      end
      test_b1_S7048: begin
        IMAGE_addr <= 7032;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 310;
        test_state <= test_b1_S7049;
      end
      test_b1_S7049: begin
        IMAGE_addr <= 7033;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7038;
        test_state <= test_b1_S7050;
      end
      test_b1_S7050: begin
        IMAGE_addr <= 7034;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 112;
        test_state <= test_b1_S7051;
      end
      test_b1_S7051: begin
        IMAGE_addr <= 7035;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S7052;
      end
      test_b1_S7052: begin
        IMAGE_addr <= 7036;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S7053;
      end
      test_b1_S7053: begin
        IMAGE_addr <= 7037;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7054;
      end
      test_b1_S7054: begin
        IMAGE_addr <= 7038;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7055;
      end
      test_b1_S7055: begin
        IMAGE_addr <= 7039;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7031;
        test_state <= test_b1_S7056;
      end
      test_b1_S7056: begin
        IMAGE_addr <= 7040;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S7057;
      end
      test_b1_S7057: begin
        IMAGE_addr <= 7041;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7052;
        test_state <= test_b1_S7058;
      end
      test_b1_S7058: begin
        IMAGE_addr <= 7042;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S7059;
      end
      test_b1_S7059: begin
        IMAGE_addr <= 7043;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S7060;
      end
      test_b1_S7060: begin
        IMAGE_addr <= 7044;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S7061;
      end
      test_b1_S7061: begin
        IMAGE_addr <= 7045;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 109;
        test_state <= test_b1_S7062;
      end
      test_b1_S7062: begin
        IMAGE_addr <= 7046;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S7063;
      end
      test_b1_S7063: begin
        IMAGE_addr <= 7047;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 110;
        test_state <= test_b1_S7064;
      end
      test_b1_S7064: begin
        IMAGE_addr <= 7048;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S7065;
      end
      test_b1_S7065: begin
        IMAGE_addr <= 7049;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S7066;
      end
      test_b1_S7066: begin
        IMAGE_addr <= 7050;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S7067;
      end
      test_b1_S7067: begin
        IMAGE_addr <= 7051;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7068;
      end
      test_b1_S7068: begin
        IMAGE_addr <= 7052;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S7069;
      end
      test_b1_S7069: begin
        IMAGE_addr <= 7053;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7070;
      end
      test_b1_S7070: begin
        IMAGE_addr <= 7054;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S7071;
      end
      test_b1_S7071: begin
        IMAGE_addr <= 7055;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7038;
        test_state <= test_b1_S7072;
      end
      test_b1_S7072: begin
        IMAGE_addr <= 7056;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S7073;
      end
      test_b1_S7073: begin
        IMAGE_addr <= 7057;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S7074;
      end
      test_b1_S7074: begin
        IMAGE_addr <= 7058;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7075;
      end
      test_b1_S7075: begin
        IMAGE_addr <= 7059;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7076;
      end
      test_b1_S7076: begin
        IMAGE_addr <= 7060;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7014;
        test_state <= test_b1_S7077;
      end
      test_b1_S7077: begin
        IMAGE_addr <= 7061;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S7078;
      end
      test_b1_S7078: begin
        IMAGE_addr <= 7062;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7069;
        test_state <= test_b1_S7079;
      end
      test_b1_S7079: begin
        IMAGE_addr <= 7063;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S7080;
      end
      test_b1_S7080: begin
        IMAGE_addr <= 7064;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S7081;
      end
      test_b1_S7081: begin
        IMAGE_addr <= 7065;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S7082;
      end
      test_b1_S7082: begin
        IMAGE_addr <= 7066;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S7083;
      end
      test_b1_S7083: begin
        IMAGE_addr <= 7067;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S7084;
      end
      test_b1_S7084: begin
        IMAGE_addr <= 7068;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7085;
      end
      test_b1_S7085: begin
        IMAGE_addr <= 7069;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7086;
      end
      test_b1_S7086: begin
        IMAGE_addr <= 7070;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7087;
      end
      test_b1_S7087: begin
        IMAGE_addr <= 7071;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S7088;
      end
      test_b1_S7088: begin
        IMAGE_addr <= 7072;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7030;
        test_state <= test_b1_S7089;
      end
      test_b1_S7089: begin
        IMAGE_addr <= 7073;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S7090;
      end
      test_b1_S7090: begin
        IMAGE_addr <= 7074;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7091;
      end
      test_b1_S7091: begin
        IMAGE_addr <= 7075;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7092;
      end
      test_b1_S7092: begin
        IMAGE_addr <= 7076;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7060;
        test_state <= test_b1_S7093;
      end
      test_b1_S7093: begin
        IMAGE_addr <= 7077;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S7094;
      end
      test_b1_S7094: begin
        IMAGE_addr <= 7078;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7083;
        test_state <= test_b1_S7095;
      end
      test_b1_S7095: begin
        IMAGE_addr <= 7079;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S7096;
      end
      test_b1_S7096: begin
        IMAGE_addr <= 7080;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 110;
        test_state <= test_b1_S7097;
      end
      test_b1_S7097: begin
        IMAGE_addr <= 7081;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 100;
        test_state <= test_b1_S7098;
      end
      test_b1_S7098: begin
        IMAGE_addr <= 7082;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7099;
      end
      test_b1_S7099: begin
        IMAGE_addr <= 7083;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7100;
      end
      test_b1_S7100: begin
        IMAGE_addr <= 7084;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7101;
      end
      test_b1_S7101: begin
        IMAGE_addr <= 7085;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S7102;
      end
      test_b1_S7102: begin
        IMAGE_addr <= 7086;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7038;
        test_state <= test_b1_S7103;
      end
      test_b1_S7103: begin
        IMAGE_addr <= 7087;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S7104;
      end
      test_b1_S7104: begin
        IMAGE_addr <= 7088;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7105;
      end
      test_b1_S7105: begin
        IMAGE_addr <= 7089;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7106;
      end
      test_b1_S7106: begin
        IMAGE_addr <= 7090;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7076;
        test_state <= test_b1_S7107;
      end
      test_b1_S7107: begin
        IMAGE_addr <= 7091;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S7108;
      end
      test_b1_S7108: begin
        IMAGE_addr <= 7092;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7097;
        test_state <= test_b1_S7109;
      end
      test_b1_S7109: begin
        IMAGE_addr <= 7093;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S7110;
      end
      test_b1_S7110: begin
        IMAGE_addr <= 7094;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 100;
        test_state <= test_b1_S7111;
      end
      test_b1_S7111: begin
        IMAGE_addr <= 7095;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 100;
        test_state <= test_b1_S7112;
      end
      test_b1_S7112: begin
        IMAGE_addr <= 7096;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7113;
      end
      test_b1_S7113: begin
        IMAGE_addr <= 7097;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7114;
      end
      test_b1_S7114: begin
        IMAGE_addr <= 7098;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7115;
      end
      test_b1_S7115: begin
        IMAGE_addr <= 7099;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7083;
        test_state <= test_b1_S7116;
      end
      test_b1_S7116: begin
        IMAGE_addr <= 7100;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S7117;
      end
      test_b1_S7117: begin
        IMAGE_addr <= 7101;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S7118;
      end
      test_b1_S7118: begin
        IMAGE_addr <= 7102;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7038;
        test_state <= test_b1_S7119;
      end
      test_b1_S7119: begin
        IMAGE_addr <= 7103;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2651;
        test_state <= test_b1_S7120;
      end
      test_b1_S7120: begin
        IMAGE_addr <= 7104;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7052;
        test_state <= test_b1_S7121;
      end
      test_b1_S7121: begin
        IMAGE_addr <= 7105;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7122;
      end
      test_b1_S7122: begin
        IMAGE_addr <= 7106;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7123;
      end
      test_b1_S7123: begin
        IMAGE_addr <= 7107;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7090;
        test_state <= test_b1_S7124;
      end
      test_b1_S7124: begin
        IMAGE_addr <= 7108;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S7125;
      end
      test_b1_S7125: begin
        IMAGE_addr <= 7109;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7114;
        test_state <= test_b1_S7126;
      end
      test_b1_S7126: begin
        IMAGE_addr <= 7110;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 103;
        test_state <= test_b1_S7127;
      end
      test_b1_S7127: begin
        IMAGE_addr <= 7111;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S7128;
      end
      test_b1_S7128: begin
        IMAGE_addr <= 7112;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S7129;
      end
      test_b1_S7129: begin
        IMAGE_addr <= 7113;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7130;
      end
      test_b1_S7130: begin
        IMAGE_addr <= 7114;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7131;
      end
      test_b1_S7131: begin
        IMAGE_addr <= 7115;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7132;
      end
      test_b1_S7132: begin
        IMAGE_addr <= 7116;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S7133;
      end
      test_b1_S7133: begin
        IMAGE_addr <= 7117;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7038;
        test_state <= test_b1_S7134;
      end
      test_b1_S7134: begin
        IMAGE_addr <= 7118;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2665;
        test_state <= test_b1_S7135;
      end
      test_b1_S7135: begin
        IMAGE_addr <= 7119;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7083;
        test_state <= test_b1_S7136;
      end
      test_b1_S7136: begin
        IMAGE_addr <= 7120;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S7137;
      end
      test_b1_S7137: begin
        IMAGE_addr <= 7121;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7052;
        test_state <= test_b1_S7138;
      end
      test_b1_S7138: begin
        IMAGE_addr <= 7122;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7139;
      end
      test_b1_S7139: begin
        IMAGE_addr <= 7123;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7140;
      end
      test_b1_S7140: begin
        IMAGE_addr <= 7124;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7107;
        test_state <= test_b1_S7141;
      end
      test_b1_S7141: begin
        IMAGE_addr <= 7125;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S7142;
      end
      test_b1_S7142: begin
        IMAGE_addr <= 7126;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7133;
        test_state <= test_b1_S7143;
      end
      test_b1_S7143: begin
        IMAGE_addr <= 7127;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S7144;
      end
      test_b1_S7144: begin
        IMAGE_addr <= 7128;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 109;
        test_state <= test_b1_S7145;
      end
      test_b1_S7145: begin
        IMAGE_addr <= 7129;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 112;
        test_state <= test_b1_S7146;
      end
      test_b1_S7146: begin
        IMAGE_addr <= 7130;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S7147;
      end
      test_b1_S7147: begin
        IMAGE_addr <= 7131;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 121;
        test_state <= test_b1_S7148;
      end
      test_b1_S7148: begin
        IMAGE_addr <= 7132;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7149;
      end
      test_b1_S7149: begin
        IMAGE_addr <= 7133;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7150;
      end
      test_b1_S7150: begin
        IMAGE_addr <= 7134;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7151;
      end
      test_b1_S7151: begin
        IMAGE_addr <= 7135;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7069;
        test_state <= test_b1_S7152;
      end
      test_b1_S7152: begin
        IMAGE_addr <= 7136;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S7153;
      end
      test_b1_S7153: begin
        IMAGE_addr <= 7137;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7038;
        test_state <= test_b1_S7154;
      end
      test_b1_S7154: begin
        IMAGE_addr <= 7138;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S7155;
      end
      test_b1_S7155: begin
        IMAGE_addr <= 7139;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7052;
        test_state <= test_b1_S7156;
      end
      test_b1_S7156: begin
        IMAGE_addr <= 7140;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7157;
      end
      test_b1_S7157: begin
        IMAGE_addr <= 7141;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7158;
      end
      test_b1_S7158: begin
        IMAGE_addr <= 7142;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7124;
        test_state <= test_b1_S7159;
      end
      test_b1_S7159: begin
        IMAGE_addr <= 7143;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S7160;
      end
      test_b1_S7160: begin
        IMAGE_addr <= 7144;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7150;
        test_state <= test_b1_S7161;
      end
      test_b1_S7161: begin
        IMAGE_addr <= 7145;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S7162;
      end
      test_b1_S7162: begin
        IMAGE_addr <= 7146;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S7163;
      end
      test_b1_S7163: begin
        IMAGE_addr <= 7147;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 122;
        test_state <= test_b1_S7164;
      end
      test_b1_S7164: begin
        IMAGE_addr <= 7148;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S7165;
      end
      test_b1_S7165: begin
        IMAGE_addr <= 7149;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7166;
      end
      test_b1_S7166: begin
        IMAGE_addr <= 7150;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7167;
      end
      test_b1_S7167: begin
        IMAGE_addr <= 7151;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7168;
      end
      test_b1_S7168: begin
        IMAGE_addr <= 7152;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7083;
        test_state <= test_b1_S7169;
      end
      test_b1_S7169: begin
        IMAGE_addr <= 7153;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7069;
        test_state <= test_b1_S7170;
      end
      test_b1_S7170: begin
        IMAGE_addr <= 7154;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 17;
        test_state <= test_b1_S7171;
      end
      test_b1_S7171: begin
        IMAGE_addr <= 7155;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7172;
      end
      test_b1_S7172: begin
        IMAGE_addr <= 7156;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7173;
      end
      test_b1_S7173: begin
        IMAGE_addr <= 7157;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7142;
        test_state <= test_b1_S7174;
      end
      test_b1_S7174: begin
        IMAGE_addr <= 7158;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S7175;
      end
      test_b1_S7175: begin
        IMAGE_addr <= 7159;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7164;
        test_state <= test_b1_S7176;
      end
      test_b1_S7176: begin
        IMAGE_addr <= 7160;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S7177;
      end
      test_b1_S7177: begin
        IMAGE_addr <= 7161;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S7178;
      end
      test_b1_S7178: begin
        IMAGE_addr <= 7162;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S7179;
      end
      test_b1_S7179: begin
        IMAGE_addr <= 7163;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7180;
      end
      test_b1_S7180: begin
        IMAGE_addr <= 7164;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7181;
      end
      test_b1_S7181: begin
        IMAGE_addr <= 7165;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7182;
      end
      test_b1_S7182: begin
        IMAGE_addr <= 7166;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S7183;
      end
      test_b1_S7183: begin
        IMAGE_addr <= 7167;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7030;
        test_state <= test_b1_S7184;
      end
      test_b1_S7184: begin
        IMAGE_addr <= 7168;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S7185;
      end
      test_b1_S7185: begin
        IMAGE_addr <= 7169;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7133;
        test_state <= test_b1_S7186;
      end
      test_b1_S7186: begin
        IMAGE_addr <= 7170;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7187;
      end
      test_b1_S7187: begin
        IMAGE_addr <= 7171;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7188;
      end
      test_b1_S7188: begin
        IMAGE_addr <= 7172;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7002;
        test_state <= test_b1_S7189;
      end
      test_b1_S7189: begin
        IMAGE_addr <= 7173;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5034;
        test_state <= test_b1_S7190;
      end
      test_b1_S7190: begin
        IMAGE_addr <= 7174;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7933;
        test_state <= test_b1_S7191;
      end
      test_b1_S7191: begin
        IMAGE_addr <= 7175;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S7192;
      end
      test_b1_S7192: begin
        IMAGE_addr <= 7176;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S7193;
      end
      test_b1_S7193: begin
        IMAGE_addr <= 7177;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S7194;
      end
      test_b1_S7194: begin
        IMAGE_addr <= 7178;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S7195;
      end
      test_b1_S7195: begin
        IMAGE_addr <= 7179;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 110;
        test_state <= test_b1_S7196;
      end
      test_b1_S7196: begin
        IMAGE_addr <= 7180;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 103;
        test_state <= test_b1_S7197;
      end
      test_b1_S7197: begin
        IMAGE_addr <= 7181;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S7198;
      end
      test_b1_S7198: begin
        IMAGE_addr <= 7182;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 39;
        test_state <= test_b1_S7199;
      end
      test_b1_S7199: begin
        IMAGE_addr <= 7183;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7200;
      end
      test_b1_S7200: begin
        IMAGE_addr <= 7184;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7201;
      end
      test_b1_S7201: begin
        IMAGE_addr <= 7185;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7202;
      end
      test_b1_S7202: begin
        IMAGE_addr <= 7186;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 306;
        test_state <= test_b1_S7203;
      end
      test_b1_S7203: begin
        IMAGE_addr <= 7187;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4956;
        test_state <= test_b1_S7204;
      end
      test_b1_S7204: begin
        IMAGE_addr <= 7188;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 37;
        test_state <= test_b1_S7205;
      end
      test_b1_S7205: begin
        IMAGE_addr <= 7189;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 37;
        test_state <= test_b1_S7206;
      end
      test_b1_S7206: begin
        IMAGE_addr <= 7190;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7207;
      end
      test_b1_S7207: begin
        IMAGE_addr <= 7191;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7185;
        test_state <= test_b1_S7208;
      end
      test_b1_S7208: begin
        IMAGE_addr <= 7192;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 310;
        test_state <= test_b1_S7209;
      end
      test_b1_S7209: begin
        IMAGE_addr <= 7193;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7198;
        test_state <= test_b1_S7210;
      end
      test_b1_S7210: begin
        IMAGE_addr <= 7194;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 108;
        test_state <= test_b1_S7211;
      end
      test_b1_S7211: begin
        IMAGE_addr <= 7195;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S7212;
      end
      test_b1_S7212: begin
        IMAGE_addr <= 7196;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 110;
        test_state <= test_b1_S7213;
      end
      test_b1_S7213: begin
        IMAGE_addr <= 7197;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7214;
      end
      test_b1_S7214: begin
        IMAGE_addr <= 7198;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7215;
      end
      test_b1_S7215: begin
        IMAGE_addr <= 7199;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7191;
        test_state <= test_b1_S7216;
      end
      test_b1_S7216: begin
        IMAGE_addr <= 7200;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 310;
        test_state <= test_b1_S7217;
      end
      test_b1_S7217: begin
        IMAGE_addr <= 7201;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7209;
        test_state <= test_b1_S7218;
      end
      test_b1_S7218: begin
        IMAGE_addr <= 7202;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 110;
        test_state <= test_b1_S7219;
      end
      test_b1_S7219: begin
        IMAGE_addr <= 7203;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S7220;
      end
      test_b1_S7220: begin
        IMAGE_addr <= 7204;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S7221;
      end
      test_b1_S7221: begin
        IMAGE_addr <= 7205;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 100;
        test_state <= test_b1_S7222;
      end
      test_b1_S7222: begin
        IMAGE_addr <= 7206;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 108;
        test_state <= test_b1_S7223;
      end
      test_b1_S7223: begin
        IMAGE_addr <= 7207;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S7224;
      end
      test_b1_S7224: begin
        IMAGE_addr <= 7208;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7225;
      end
      test_b1_S7225: begin
        IMAGE_addr <= 7209;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7226;
      end
      test_b1_S7226: begin
        IMAGE_addr <= 7210;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7199;
        test_state <= test_b1_S7227;
      end
      test_b1_S7227: begin
        IMAGE_addr <= 7211;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 310;
        test_state <= test_b1_S7228;
      end
      test_b1_S7228: begin
        IMAGE_addr <= 7212;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7222;
        test_state <= test_b1_S7229;
      end
      test_b1_S7229: begin
        IMAGE_addr <= 7213;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 104;
        test_state <= test_b1_S7230;
      end
      test_b1_S7230: begin
        IMAGE_addr <= 7214;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S7231;
      end
      test_b1_S7231: begin
        IMAGE_addr <= 7215;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 121;
        test_state <= test_b1_S7232;
      end
      test_b1_S7232: begin
        IMAGE_addr <= 7216;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S7233;
      end
      test_b1_S7233: begin
        IMAGE_addr <= 7217;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S7234;
      end
      test_b1_S7234: begin
        IMAGE_addr <= 7218;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S7235;
      end
      test_b1_S7235: begin
        IMAGE_addr <= 7219;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 99;
        test_state <= test_b1_S7236;
      end
      test_b1_S7236: begin
        IMAGE_addr <= 7220;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 107;
        test_state <= test_b1_S7237;
      end
      test_b1_S7237: begin
        IMAGE_addr <= 7221;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7238;
      end
      test_b1_S7238: begin
        IMAGE_addr <= 7222;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7239;
      end
      test_b1_S7239: begin
        IMAGE_addr <= 7223;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7210;
        test_state <= test_b1_S7240;
      end
      test_b1_S7240: begin
        IMAGE_addr <= 7224;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 310;
        test_state <= test_b1_S7241;
      end
      test_b1_S7241: begin
        IMAGE_addr <= 7225;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7231;
        test_state <= test_b1_S7242;
      end
      test_b1_S7242: begin
        IMAGE_addr <= 7226;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 102;
        test_state <= test_b1_S7243;
      end
      test_b1_S7243: begin
        IMAGE_addr <= 7227;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 108;
        test_state <= test_b1_S7244;
      end
      test_b1_S7244: begin
        IMAGE_addr <= 7228;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S7245;
      end
      test_b1_S7245: begin
        IMAGE_addr <= 7229;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 103;
        test_state <= test_b1_S7246;
      end
      test_b1_S7246: begin
        IMAGE_addr <= 7230;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7247;
      end
      test_b1_S7247: begin
        IMAGE_addr <= 7231;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7248;
      end
      test_b1_S7248: begin
        IMAGE_addr <= 7232;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7223;
        test_state <= test_b1_S7249;
      end
      test_b1_S7249: begin
        IMAGE_addr <= 7233;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 310;
        test_state <= test_b1_S7250;
      end
      test_b1_S7250: begin
        IMAGE_addr <= 7234;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7241;
        test_state <= test_b1_S7251;
      end
      test_b1_S7251: begin
        IMAGE_addr <= 7235;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S7252;
      end
      test_b1_S7252: begin
        IMAGE_addr <= 7236;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S7253;
      end
      test_b1_S7253: begin
        IMAGE_addr <= 7237;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 103;
        test_state <= test_b1_S7254;
      end
      test_b1_S7254: begin
        IMAGE_addr <= 7238;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 104;
        test_state <= test_b1_S7255;
      end
      test_b1_S7255: begin
        IMAGE_addr <= 7239;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S7256;
      end
      test_b1_S7256: begin
        IMAGE_addr <= 7240;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7257;
      end
      test_b1_S7257: begin
        IMAGE_addr <= 7241;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7258;
      end
      test_b1_S7258: begin
        IMAGE_addr <= 7242;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7232;
        test_state <= test_b1_S7259;
      end
      test_b1_S7259: begin
        IMAGE_addr <= 7243;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 310;
        test_state <= test_b1_S7260;
      end
      test_b1_S7260: begin
        IMAGE_addr <= 7244;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7250;
        test_state <= test_b1_S7261;
      end
      test_b1_S7261: begin
        IMAGE_addr <= 7245;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 108;
        test_state <= test_b1_S7262;
      end
      test_b1_S7262: begin
        IMAGE_addr <= 7246;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S7263;
      end
      test_b1_S7263: begin
        IMAGE_addr <= 7247;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 102;
        test_state <= test_b1_S7264;
      end
      test_b1_S7264: begin
        IMAGE_addr <= 7248;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S7265;
      end
      test_b1_S7265: begin
        IMAGE_addr <= 7249;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7266;
      end
      test_b1_S7266: begin
        IMAGE_addr <= 7250;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7267;
      end
      test_b1_S7267: begin
        IMAGE_addr <= 7251;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7242;
        test_state <= test_b1_S7268;
      end
      test_b1_S7268: begin
        IMAGE_addr <= 7252;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 310;
        test_state <= test_b1_S7269;
      end
      test_b1_S7269: begin
        IMAGE_addr <= 7253;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7258;
        test_state <= test_b1_S7270;
      end
      test_b1_S7270: begin
        IMAGE_addr <= 7254;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S7271;
      end
      test_b1_S7271: begin
        IMAGE_addr <= 7255;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S7272;
      end
      test_b1_S7272: begin
        IMAGE_addr <= 7256;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 99;
        test_state <= test_b1_S7273;
      end
      test_b1_S7273: begin
        IMAGE_addr <= 7257;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7274;
      end
      test_b1_S7274: begin
        IMAGE_addr <= 7258;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7275;
      end
      test_b1_S7275: begin
        IMAGE_addr <= 7259;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7251;
        test_state <= test_b1_S7276;
      end
      test_b1_S7276: begin
        IMAGE_addr <= 7260;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S7277;
      end
      test_b1_S7277: begin
        IMAGE_addr <= 7261;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7269;
        test_state <= test_b1_S7278;
      end
      test_b1_S7278: begin
        IMAGE_addr <= 7262;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 98;
        test_state <= test_b1_S7279;
      end
      test_b1_S7279: begin
        IMAGE_addr <= 7263;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 117;
        test_state <= test_b1_S7280;
      end
      test_b1_S7280: begin
        IMAGE_addr <= 7264;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 102;
        test_state <= test_b1_S7281;
      end
      test_b1_S7281: begin
        IMAGE_addr <= 7265;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 102;
        test_state <= test_b1_S7282;
      end
      test_b1_S7282: begin
        IMAGE_addr <= 7266;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S7283;
      end
      test_b1_S7283: begin
        IMAGE_addr <= 7267;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S7284;
      end
      test_b1_S7284: begin
        IMAGE_addr <= 7268;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7285;
      end
      test_b1_S7285: begin
        IMAGE_addr <= 7269;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 206;
        test_state <= test_b1_S7286;
      end
      test_b1_S7286: begin
        IMAGE_addr <= 7270;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 909;
        test_state <= test_b1_S7287;
      end
      test_b1_S7287: begin
        IMAGE_addr <= 7271;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S7288;
      end
      test_b1_S7288: begin
        IMAGE_addr <= 7272;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S7289;
      end
      test_b1_S7289: begin
        IMAGE_addr <= 7273;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 18;
        test_state <= test_b1_S7290;
      end
      test_b1_S7290: begin
        IMAGE_addr <= 7274;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 16;
        test_state <= test_b1_S7291;
      end
      test_b1_S7291: begin
        IMAGE_addr <= 7275;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 915;
        test_state <= test_b1_S7292;
      end
      test_b1_S7292: begin
        IMAGE_addr <= 7276;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 909;
        test_state <= test_b1_S7293;
      end
      test_b1_S7293: begin
        IMAGE_addr <= 7277;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 18;
        test_state <= test_b1_S7294;
      end
      test_b1_S7294: begin
        IMAGE_addr <= 7278;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 16;
        test_state <= test_b1_S7295;
      end
      test_b1_S7295: begin
        IMAGE_addr <= 7279;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7296;
      end
      test_b1_S7296: begin
        IMAGE_addr <= 7280;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7297;
      end
      test_b1_S7297: begin
        IMAGE_addr <= 7281;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7259;
        test_state <= test_b1_S7298;
      end
      test_b1_S7298: begin
        IMAGE_addr <= 7282;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S7299;
      end
      test_b1_S7299: begin
        IMAGE_addr <= 7283;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7289;
        test_state <= test_b1_S7300;
      end
      test_b1_S7300: begin
        IMAGE_addr <= 7284;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S7301;
      end
      test_b1_S7301: begin
        IMAGE_addr <= 7285;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S7302;
      end
      test_b1_S7302: begin
        IMAGE_addr <= 7286;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S7303;
      end
      test_b1_S7303: begin
        IMAGE_addr <= 7287;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 109;
        test_state <= test_b1_S7304;
      end
      test_b1_S7304: begin
        IMAGE_addr <= 7288;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7305;
      end
      test_b1_S7305: begin
        IMAGE_addr <= 7289;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S7306;
      end
      test_b1_S7306: begin
        IMAGE_addr <= 7290;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 886;
        test_state <= test_b1_S7307;
      end
      test_b1_S7307: begin
        IMAGE_addr <= 7291;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 16;
        test_state <= test_b1_S7308;
      end
      test_b1_S7308: begin
        IMAGE_addr <= 7292;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 27;
        test_state <= test_b1_S7309;
      end
      test_b1_S7309: begin
        IMAGE_addr <= 7293;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S7310;
      end
      test_b1_S7310: begin
        IMAGE_addr <= 7294;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S7311;
      end
      test_b1_S7311: begin
        IMAGE_addr <= 7295;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S7312;
      end
      test_b1_S7312: begin
        IMAGE_addr <= 7296;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 32;
        test_state <= test_b1_S7313;
      end
      test_b1_S7313: begin
        IMAGE_addr <= 7297;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 790;
        test_state <= test_b1_S7314;
      end
      test_b1_S7314: begin
        IMAGE_addr <= 7298;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S7315;
      end
      test_b1_S7315: begin
        IMAGE_addr <= 7299;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7309;
        test_state <= test_b1_S7316;
      end
      test_b1_S7316: begin
        IMAGE_addr <= 7300;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S7317;
      end
      test_b1_S7317: begin
        IMAGE_addr <= 7301;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7318;
      end
      test_b1_S7318: begin
        IMAGE_addr <= 7302;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S7319;
      end
      test_b1_S7319: begin
        IMAGE_addr <= 7303;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S7320;
      end
      test_b1_S7320: begin
        IMAGE_addr <= 7304;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S7321;
      end
      test_b1_S7321: begin
        IMAGE_addr <= 7305;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 27;
        test_state <= test_b1_S7322;
      end
      test_b1_S7322: begin
        IMAGE_addr <= 7306;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2665;
        test_state <= test_b1_S7323;
      end
      test_b1_S7323: begin
        IMAGE_addr <= 7307;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7289;
        test_state <= test_b1_S7324;
      end
      test_b1_S7324: begin
        IMAGE_addr <= 7308;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7325;
      end
      test_b1_S7325: begin
        IMAGE_addr <= 7309;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S7326;
      end
      test_b1_S7326: begin
        IMAGE_addr <= 7310;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 52;
        test_state <= test_b1_S7327;
      end
      test_b1_S7327: begin
        IMAGE_addr <= 7311;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 732;
        test_state <= test_b1_S7328;
      end
      test_b1_S7328: begin
        IMAGE_addr <= 7312;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7329;
      end
      test_b1_S7329: begin
        IMAGE_addr <= 7313;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7330;
      end
      test_b1_S7330: begin
        IMAGE_addr <= 7314;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7281;
        test_state <= test_b1_S7331;
      end
      test_b1_S7331: begin
        IMAGE_addr <= 7315;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S7332;
      end
      test_b1_S7332: begin
        IMAGE_addr <= 7316;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7323;
        test_state <= test_b1_S7333;
      end
      test_b1_S7333: begin
        IMAGE_addr <= 7317;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 112;
        test_state <= test_b1_S7334;
      end
      test_b1_S7334: begin
        IMAGE_addr <= 7318;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 108;
        test_state <= test_b1_S7335;
      end
      test_b1_S7335: begin
        IMAGE_addr <= 7319;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S7336;
      end
      test_b1_S7336: begin
        IMAGE_addr <= 7320;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 99;
        test_state <= test_b1_S7337;
      end
      test_b1_S7337: begin
        IMAGE_addr <= 7321;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S7338;
      end
      test_b1_S7338: begin
        IMAGE_addr <= 7322;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7339;
      end
      test_b1_S7339: begin
        IMAGE_addr <= 7323;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S7340;
      end
      test_b1_S7340: begin
        IMAGE_addr <= 7324;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7329;
        test_state <= test_b1_S7341;
      end
      test_b1_S7341: begin
        IMAGE_addr <= 7325;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4126;
        test_state <= test_b1_S7342;
      end
      test_b1_S7342: begin
        IMAGE_addr <= 7326;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S7343;
      end
      test_b1_S7343: begin
        IMAGE_addr <= 7327;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7344;
      end
      test_b1_S7344: begin
        IMAGE_addr <= 7328;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7345;
      end
      test_b1_S7345: begin
        IMAGE_addr <= 7329;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 774;
        test_state <= test_b1_S7346;
      end
      test_b1_S7346: begin
        IMAGE_addr <= 7330;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 206;
        test_state <= test_b1_S7347;
      end
      test_b1_S7347: begin
        IMAGE_addr <= 7331;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 16;
        test_state <= test_b1_S7348;
      end
      test_b1_S7348: begin
        IMAGE_addr <= 7332;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S7349;
      end
      test_b1_S7349: begin
        IMAGE_addr <= 7333;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7350;
      end
      test_b1_S7350: begin
        IMAGE_addr <= 7334;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7351;
      end
      test_b1_S7351: begin
        IMAGE_addr <= 7335;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7314;
        test_state <= test_b1_S7352;
      end
      test_b1_S7352: begin
        IMAGE_addr <= 7336;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S7353;
      end
      test_b1_S7353: begin
        IMAGE_addr <= 7337;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7343;
        test_state <= test_b1_S7354;
      end
      test_b1_S7354: begin
        IMAGE_addr <= 7338;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 112;
        test_state <= test_b1_S7355;
      end
      test_b1_S7355: begin
        IMAGE_addr <= 7339;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S7356;
      end
      test_b1_S7356: begin
        IMAGE_addr <= 7340;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S7357;
      end
      test_b1_S7357: begin
        IMAGE_addr <= 7341;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 112;
        test_state <= test_b1_S7358;
      end
      test_b1_S7358: begin
        IMAGE_addr <= 7342;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7359;
      end
      test_b1_S7359: begin
        IMAGE_addr <= 7343;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S7360;
      end
      test_b1_S7360: begin
        IMAGE_addr <= 7344;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S7361;
      end
      test_b1_S7361: begin
        IMAGE_addr <= 7345;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7222;
        test_state <= test_b1_S7362;
      end
      test_b1_S7362: begin
        IMAGE_addr <= 7346;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S7363;
      end
      test_b1_S7363: begin
        IMAGE_addr <= 7347;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S7364;
      end
      test_b1_S7364: begin
        IMAGE_addr <= 7348;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7354;
        test_state <= test_b1_S7365;
      end
      test_b1_S7365: begin
        IMAGE_addr <= 7349;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 877;
        test_state <= test_b1_S7366;
      end
      test_b1_S7366: begin
        IMAGE_addr <= 7350;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S7367;
      end
      test_b1_S7367: begin
        IMAGE_addr <= 7351;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7198;
        test_state <= test_b1_S7368;
      end
      test_b1_S7368: begin
        IMAGE_addr <= 7352;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S7369;
      end
      test_b1_S7369: begin
        IMAGE_addr <= 7353;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7370;
      end
      test_b1_S7370: begin
        IMAGE_addr <= 7354;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S7371;
      end
      test_b1_S7371: begin
        IMAGE_addr <= 7355;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7360;
        test_state <= test_b1_S7372;
      end
      test_b1_S7372: begin
        IMAGE_addr <= 7356;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S7373;
      end
      test_b1_S7373: begin
        IMAGE_addr <= 7357;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7209;
        test_state <= test_b1_S7374;
      end
      test_b1_S7374: begin
        IMAGE_addr <= 7358;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S7375;
      end
      test_b1_S7375: begin
        IMAGE_addr <= 7359;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7376;
      end
      test_b1_S7376: begin
        IMAGE_addr <= 7360;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3539;
        test_state <= test_b1_S7377;
      end
      test_b1_S7377: begin
        IMAGE_addr <= 7361;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S7378;
      end
      test_b1_S7378: begin
        IMAGE_addr <= 7362;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7379;
      end
      test_b1_S7379: begin
        IMAGE_addr <= 7363;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S7380;
      end
      test_b1_S7380: begin
        IMAGE_addr <= 7364;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7231;
        test_state <= test_b1_S7381;
      end
      test_b1_S7381: begin
        IMAGE_addr <= 7365;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S7382;
      end
      test_b1_S7382: begin
        IMAGE_addr <= 7366;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7383;
      end
      test_b1_S7383: begin
        IMAGE_addr <= 7367;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7384;
      end
      test_b1_S7384: begin
        IMAGE_addr <= 7368;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7335;
        test_state <= test_b1_S7385;
      end
      test_b1_S7385: begin
        IMAGE_addr <= 7369;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S7386;
      end
      test_b1_S7386: begin
        IMAGE_addr <= 7370;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7376;
        test_state <= test_b1_S7387;
      end
      test_b1_S7387: begin
        IMAGE_addr <= 7371;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 109;
        test_state <= test_b1_S7388;
      end
      test_b1_S7388: begin
        IMAGE_addr <= 7372;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 111;
        test_state <= test_b1_S7389;
      end
      test_b1_S7389: begin
        IMAGE_addr <= 7373;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 118;
        test_state <= test_b1_S7390;
      end
      test_b1_S7390: begin
        IMAGE_addr <= 7374;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S7391;
      end
      test_b1_S7391: begin
        IMAGE_addr <= 7375;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7392;
      end
      test_b1_S7392: begin
        IMAGE_addr <= 7376;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S7393;
      end
      test_b1_S7393: begin
        IMAGE_addr <= 7377;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7222;
        test_state <= test_b1_S7394;
      end
      test_b1_S7394: begin
        IMAGE_addr <= 7378;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S7395;
      end
      test_b1_S7395: begin
        IMAGE_addr <= 7379;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 206;
        test_state <= test_b1_S7396;
      end
      test_b1_S7396: begin
        IMAGE_addr <= 7380;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S7397;
      end
      test_b1_S7397: begin
        IMAGE_addr <= 7381;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7198;
        test_state <= test_b1_S7398;
      end
      test_b1_S7398: begin
        IMAGE_addr <= 7382;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S7399;
      end
      test_b1_S7399: begin
        IMAGE_addr <= 7383;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7323;
        test_state <= test_b1_S7400;
      end
      test_b1_S7400: begin
        IMAGE_addr <= 7384;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S7401;
      end
      test_b1_S7401: begin
        IMAGE_addr <= 7385;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7222;
        test_state <= test_b1_S7402;
      end
      test_b1_S7402: begin
        IMAGE_addr <= 7386;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2651;
        test_state <= test_b1_S7403;
      end
      test_b1_S7403: begin
        IMAGE_addr <= 7387;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7404;
      end
      test_b1_S7404: begin
        IMAGE_addr <= 7388;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7405;
      end
      test_b1_S7405: begin
        IMAGE_addr <= 7389;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7368;
        test_state <= test_b1_S7406;
      end
      test_b1_S7406: begin
        IMAGE_addr <= 7390;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S7407;
      end
      test_b1_S7407: begin
        IMAGE_addr <= 7391;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7396;
        test_state <= test_b1_S7408;
      end
      test_b1_S7408: begin
        IMAGE_addr <= 7392;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 99;
        test_state <= test_b1_S7409;
      end
      test_b1_S7409: begin
        IMAGE_addr <= 7393;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 109;
        test_state <= test_b1_S7410;
      end
      test_b1_S7410: begin
        IMAGE_addr <= 7394;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 112;
        test_state <= test_b1_S7411;
      end
      test_b1_S7411: begin
        IMAGE_addr <= 7395;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7412;
      end
      test_b1_S7412: begin
        IMAGE_addr <= 7396;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S7413;
      end
      test_b1_S7413: begin
        IMAGE_addr <= 7397;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7231;
        test_state <= test_b1_S7414;
      end
      test_b1_S7414: begin
        IMAGE_addr <= 7398;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S7415;
      end
      test_b1_S7415: begin
        IMAGE_addr <= 7399;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S7416;
      end
      test_b1_S7416: begin
        IMAGE_addr <= 7400;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7417;
      end
      test_b1_S7417: begin
        IMAGE_addr <= 7401;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 798;
        test_state <= test_b1_S7418;
      end
      test_b1_S7418: begin
        IMAGE_addr <= 7402;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 140;
        test_state <= test_b1_S7419;
      end
      test_b1_S7419: begin
        IMAGE_addr <= 7403;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 25;
        test_state <= test_b1_S7420;
      end
      test_b1_S7420: begin
        IMAGE_addr <= 7404;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S7421;
      end
      test_b1_S7421: begin
        IMAGE_addr <= 7405;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S7422;
      end
      test_b1_S7422: begin
        IMAGE_addr <= 7406;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7209;
        test_state <= test_b1_S7423;
      end
      test_b1_S7423: begin
        IMAGE_addr <= 7407;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S7424;
      end
      test_b1_S7424: begin
        IMAGE_addr <= 7408;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 206;
        test_state <= test_b1_S7425;
      end
      test_b1_S7425: begin
        IMAGE_addr <= 7409;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 838;
        test_state <= test_b1_S7426;
      end
      test_b1_S7426: begin
        IMAGE_addr <= 7410;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S7427;
      end
      test_b1_S7427: begin
        IMAGE_addr <= 7411;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7420;
        test_state <= test_b1_S7428;
      end
      test_b1_S7428: begin
        IMAGE_addr <= 7412;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S7429;
      end
      test_b1_S7429: begin
        IMAGE_addr <= 7413;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7222;
        test_state <= test_b1_S7430;
      end
      test_b1_S7430: begin
        IMAGE_addr <= 7414;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S7431;
      end
      test_b1_S7431: begin
        IMAGE_addr <= 7415;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 27;
        test_state <= test_b1_S7432;
      end
      test_b1_S7432: begin
        IMAGE_addr <= 7416;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S7433;
      end
      test_b1_S7433: begin
        IMAGE_addr <= 7417;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7231;
        test_state <= test_b1_S7434;
      end
      test_b1_S7434: begin
        IMAGE_addr <= 7418;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S7435;
      end
      test_b1_S7435: begin
        IMAGE_addr <= 7419;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7436;
      end
      test_b1_S7436: begin
        IMAGE_addr <= 7420;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 751;
        test_state <= test_b1_S7437;
      end
      test_b1_S7437: begin
        IMAGE_addr <= 7421;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7438;
      end
      test_b1_S7438: begin
        IMAGE_addr <= 7422;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7439;
      end
      test_b1_S7439: begin
        IMAGE_addr <= 7423;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7185;
        test_state <= test_b1_S7440;
      end
      test_b1_S7440: begin
        IMAGE_addr <= 7424;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S7441;
      end
      test_b1_S7441: begin
        IMAGE_addr <= 7425;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7433;
        test_state <= test_b1_S7442;
      end
      test_b1_S7442: begin
        IMAGE_addr <= 7426;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S7443;
      end
      test_b1_S7443: begin
        IMAGE_addr <= 7427;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S7444;
      end
      test_b1_S7444: begin
        IMAGE_addr <= 7428;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S7445;
      end
      test_b1_S7445: begin
        IMAGE_addr <= 7429;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S7446;
      end
      test_b1_S7446: begin
        IMAGE_addr <= 7430;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 99;
        test_state <= test_b1_S7447;
      end
      test_b1_S7447: begin
        IMAGE_addr <= 7431;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 104;
        test_state <= test_b1_S7448;
      end
      test_b1_S7448: begin
        IMAGE_addr <= 7432;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7449;
      end
      test_b1_S7449: begin
        IMAGE_addr <= 7433;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7450;
      end
      test_b1_S7450: begin
        IMAGE_addr <= 7434;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7451;
      end
      test_b1_S7451: begin
        IMAGE_addr <= 7435;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S7452;
      end
      test_b1_S7452: begin
        IMAGE_addr <= 7436;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7231;
        test_state <= test_b1_S7453;
      end
      test_b1_S7453: begin
        IMAGE_addr <= 7437;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 155;
        test_state <= test_b1_S7454;
      end
      test_b1_S7454: begin
        IMAGE_addr <= 7438;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7343;
        test_state <= test_b1_S7455;
      end
      test_b1_S7455: begin
        IMAGE_addr <= 7439;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S7456;
      end
      test_b1_S7456: begin
        IMAGE_addr <= 7440;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7222;
        test_state <= test_b1_S7457;
      end
      test_b1_S7457: begin
        IMAGE_addr <= 7441;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S7458;
      end
      test_b1_S7458: begin
        IMAGE_addr <= 7442;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 877;
        test_state <= test_b1_S7459;
      end
      test_b1_S7459: begin
        IMAGE_addr <= 7443;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S7460;
      end
      test_b1_S7460: begin
        IMAGE_addr <= 7444;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7448;
        test_state <= test_b1_S7461;
      end
      test_b1_S7461: begin
        IMAGE_addr <= 7445;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7376;
        test_state <= test_b1_S7462;
      end
      test_b1_S7462: begin
        IMAGE_addr <= 7446;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7396;
        test_state <= test_b1_S7463;
      end
      test_b1_S7463: begin
        IMAGE_addr <= 7447;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7464;
      end
      test_b1_S7464: begin
        IMAGE_addr <= 7448;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3841;
        test_state <= test_b1_S7465;
      end
      test_b1_S7465: begin
        IMAGE_addr <= 7449;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S7466;
      end
      test_b1_S7466: begin
        IMAGE_addr <= 7450;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7231;
        test_state <= test_b1_S7467;
      end
      test_b1_S7467: begin
        IMAGE_addr <= 7451;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S7468;
      end
      test_b1_S7468: begin
        IMAGE_addr <= 7452;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7469;
      end
      test_b1_S7469: begin
        IMAGE_addr <= 7453;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7470;
      end
      test_b1_S7470: begin
        IMAGE_addr <= 7454;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7423;
        test_state <= test_b1_S7471;
      end
      test_b1_S7471: begin
        IMAGE_addr <= 7455;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S7472;
      end
      test_b1_S7472: begin
        IMAGE_addr <= 7456;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7466;
        test_state <= test_b1_S7473;
      end
      test_b1_S7473: begin
        IMAGE_addr <= 7457;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 102;
        test_state <= test_b1_S7474;
      end
      test_b1_S7474: begin
        IMAGE_addr <= 7458;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S7475;
      end
      test_b1_S7475: begin
        IMAGE_addr <= 7459;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 110;
        test_state <= test_b1_S7476;
      end
      test_b1_S7476: begin
        IMAGE_addr <= 7460;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 100;
        test_state <= test_b1_S7477;
      end
      test_b1_S7477: begin
        IMAGE_addr <= 7461;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 67;
        test_state <= test_b1_S7478;
      end
      test_b1_S7478: begin
        IMAGE_addr <= 7462;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 104;
        test_state <= test_b1_S7479;
      end
      test_b1_S7479: begin
        IMAGE_addr <= 7463;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S7480;
      end
      test_b1_S7480: begin
        IMAGE_addr <= 7464;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S7481;
      end
      test_b1_S7481: begin
        IMAGE_addr <= 7465;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7482;
      end
      test_b1_S7482: begin
        IMAGE_addr <= 7466;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7483;
      end
      test_b1_S7483: begin
        IMAGE_addr <= 7467;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7484;
      end
      test_b1_S7484: begin
        IMAGE_addr <= 7468;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S7485;
      end
      test_b1_S7485: begin
        IMAGE_addr <= 7469;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7209;
        test_state <= test_b1_S7486;
      end
      test_b1_S7486: begin
        IMAGE_addr <= 7470;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S7487;
      end
      test_b1_S7487: begin
        IMAGE_addr <= 7471;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 189;
        test_state <= test_b1_S7488;
      end
      test_b1_S7488: begin
        IMAGE_addr <= 7472;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S7489;
      end
      test_b1_S7489: begin
        IMAGE_addr <= 7473;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S7490;
      end
      test_b1_S7490: begin
        IMAGE_addr <= 7474;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7491;
      end
      test_b1_S7491: begin
        IMAGE_addr <= 7475;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 790;
        test_state <= test_b1_S7492;
      end
      test_b1_S7492: begin
        IMAGE_addr <= 7476;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S7493;
      end
      test_b1_S7493: begin
        IMAGE_addr <= 7477;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7485;
        test_state <= test_b1_S7494;
      end
      test_b1_S7494: begin
        IMAGE_addr <= 7478;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S7495;
      end
      test_b1_S7495: begin
        IMAGE_addr <= 7479;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S7496;
      end
      test_b1_S7496: begin
        IMAGE_addr <= 7480;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S7497;
      end
      test_b1_S7497: begin
        IMAGE_addr <= 7481;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7498;
      end
      test_b1_S7498: begin
        IMAGE_addr <= 7482;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S7499;
      end
      test_b1_S7499: begin
        IMAGE_addr <= 7483;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7500;
      end
      test_b1_S7500: begin
        IMAGE_addr <= 7484;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7501;
      end
      test_b1_S7501: begin
        IMAGE_addr <= 7485;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S7502;
      end
      test_b1_S7502: begin
        IMAGE_addr <= 7486;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7490;
        test_state <= test_b1_S7503;
      end
      test_b1_S7503: begin
        IMAGE_addr <= 7487;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S7504;
      end
      test_b1_S7504: begin
        IMAGE_addr <= 7488;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4294967295;
        test_state <= test_b1_S7505;
      end
      test_b1_S7505: begin
        IMAGE_addr <= 7489;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7506;
      end
      test_b1_S7506: begin
        IMAGE_addr <= 7490;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 732;
        test_state <= test_b1_S7507;
      end
      test_b1_S7507: begin
        IMAGE_addr <= 7491;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 25;
        test_state <= test_b1_S7508;
      end
      test_b1_S7508: begin
        IMAGE_addr <= 7492;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S7509;
      end
      test_b1_S7509: begin
        IMAGE_addr <= 7493;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S7510;
      end
      test_b1_S7510: begin
        IMAGE_addr <= 7494;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7209;
        test_state <= test_b1_S7511;
      end
      test_b1_S7511: begin
        IMAGE_addr <= 7495;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S7512;
      end
      test_b1_S7512: begin
        IMAGE_addr <= 7496;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 790;
        test_state <= test_b1_S7513;
      end
      test_b1_S7513: begin
        IMAGE_addr <= 7497;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S7514;
      end
      test_b1_S7514: begin
        IMAGE_addr <= 7498;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7503;
        test_state <= test_b1_S7515;
      end
      test_b1_S7515: begin
        IMAGE_addr <= 7499;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 27;
        test_state <= test_b1_S7516;
      end
      test_b1_S7516: begin
        IMAGE_addr <= 7500;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S7517;
      end
      test_b1_S7517: begin
        IMAGE_addr <= 7501;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7518;
      end
      test_b1_S7518: begin
        IMAGE_addr <= 7502;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7519;
      end
      test_b1_S7519: begin
        IMAGE_addr <= 7503;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S7520;
      end
      test_b1_S7520: begin
        IMAGE_addr <= 7504;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7508;
        test_state <= test_b1_S7521;
      end
      test_b1_S7521: begin
        IMAGE_addr <= 7505;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S7522;
      end
      test_b1_S7522: begin
        IMAGE_addr <= 7506;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4294967295;
        test_state <= test_b1_S7523;
      end
      test_b1_S7523: begin
        IMAGE_addr <= 7507;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7524;
      end
      test_b1_S7524: begin
        IMAGE_addr <= 7508;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 732;
        test_state <= test_b1_S7525;
      end
      test_b1_S7525: begin
        IMAGE_addr <= 7509;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 25;
        test_state <= test_b1_S7526;
      end
      test_b1_S7526: begin
        IMAGE_addr <= 7510;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S7527;
      end
      test_b1_S7527: begin
        IMAGE_addr <= 7511;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8;
        test_state <= test_b1_S7528;
      end
      test_b1_S7528: begin
        IMAGE_addr <= 7512;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7471;
        test_state <= test_b1_S7529;
      end
      test_b1_S7529: begin
        IMAGE_addr <= 7513;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7530;
      end
      test_b1_S7530: begin
        IMAGE_addr <= 7514;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7531;
      end
      test_b1_S7531: begin
        IMAGE_addr <= 7515;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7454;
        test_state <= test_b1_S7532;
      end
      test_b1_S7532: begin
        IMAGE_addr <= 7516;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S7533;
      end
      test_b1_S7533: begin
        IMAGE_addr <= 7517;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7523;
        test_state <= test_b1_S7534;
      end
      test_b1_S7534: begin
        IMAGE_addr <= 7518;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 99;
        test_state <= test_b1_S7535;
      end
      test_b1_S7535: begin
        IMAGE_addr <= 7519;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 104;
        test_state <= test_b1_S7536;
      end
      test_b1_S7536: begin
        IMAGE_addr <= 7520;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 111;
        test_state <= test_b1_S7537;
      end
      test_b1_S7537: begin
        IMAGE_addr <= 7521;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 112;
        test_state <= test_b1_S7538;
      end
      test_b1_S7538: begin
        IMAGE_addr <= 7522;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7539;
      end
      test_b1_S7539: begin
        IMAGE_addr <= 7523;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7540;
      end
      test_b1_S7540: begin
        IMAGE_addr <= 7524;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7541;
      end
      test_b1_S7541: begin
        IMAGE_addr <= 7525;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5792;
        test_state <= test_b1_S7542;
      end
      test_b1_S7542: begin
        IMAGE_addr <= 7526;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 886;
        test_state <= test_b1_S7543;
      end
      test_b1_S7543: begin
        IMAGE_addr <= 7527;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 132;
        test_state <= test_b1_S7544;
      end
      test_b1_S7544: begin
        IMAGE_addr <= 7528;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 16;
        test_state <= test_b1_S7545;
      end
      test_b1_S7545: begin
        IMAGE_addr <= 7529;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 27;
        test_state <= test_b1_S7546;
      end
      test_b1_S7546: begin
        IMAGE_addr <= 7530;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S7547;
      end
      test_b1_S7547: begin
        IMAGE_addr <= 7531;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7548;
      end
      test_b1_S7548: begin
        IMAGE_addr <= 7532;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S7549;
      end
      test_b1_S7549: begin
        IMAGE_addr <= 7533;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S7550;
      end
      test_b1_S7550: begin
        IMAGE_addr <= 7534;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7551;
      end
      test_b1_S7551: begin
        IMAGE_addr <= 7535;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7552;
      end
      test_b1_S7552: begin
        IMAGE_addr <= 7536;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7515;
        test_state <= test_b1_S7553;
      end
      test_b1_S7553: begin
        IMAGE_addr <= 7537;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S7554;
      end
      test_b1_S7554: begin
        IMAGE_addr <= 7538;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7549;
        test_state <= test_b1_S7555;
      end
      test_b1_S7555: begin
        IMAGE_addr <= 7539;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 103;
        test_state <= test_b1_S7556;
      end
      test_b1_S7556: begin
        IMAGE_addr <= 7540;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S7557;
      end
      test_b1_S7557: begin
        IMAGE_addr <= 7541;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S7558;
      end
      test_b1_S7558: begin
        IMAGE_addr <= 7542;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 83;
        test_state <= test_b1_S7559;
      end
      test_b1_S7559: begin
        IMAGE_addr <= 7543;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 117;
        test_state <= test_b1_S7560;
      end
      test_b1_S7560: begin
        IMAGE_addr <= 7544;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 98;
        test_state <= test_b1_S7561;
      end
      test_b1_S7561: begin
        IMAGE_addr <= 7545;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S7562;
      end
      test_b1_S7562: begin
        IMAGE_addr <= 7546;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S7563;
      end
      test_b1_S7563: begin
        IMAGE_addr <= 7547;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S7564;
      end
      test_b1_S7564: begin
        IMAGE_addr <= 7548;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7565;
      end
      test_b1_S7565: begin
        IMAGE_addr <= 7549;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7566;
      end
      test_b1_S7566: begin
        IMAGE_addr <= 7550;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7567;
      end
      test_b1_S7567: begin
        IMAGE_addr <= 7551;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7269;
        test_state <= test_b1_S7568;
      end
      test_b1_S7568: begin
        IMAGE_addr <= 7552;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S7569;
      end
      test_b1_S7569: begin
        IMAGE_addr <= 7553;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7570;
      end
      test_b1_S7570: begin
        IMAGE_addr <= 7554;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 909;
        test_state <= test_b1_S7571;
      end
      test_b1_S7571: begin
        IMAGE_addr <= 7555;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4148;
        test_state <= test_b1_S7572;
      end
      test_b1_S7572: begin
        IMAGE_addr <= 7556;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S7573;
      end
      test_b1_S7573: begin
        IMAGE_addr <= 7557;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7241;
        test_state <= test_b1_S7574;
      end
      test_b1_S7574: begin
        IMAGE_addr <= 7558;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S7575;
      end
      test_b1_S7575: begin
        IMAGE_addr <= 7559;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S7576;
      end
      test_b1_S7576: begin
        IMAGE_addr <= 7560;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7250;
        test_state <= test_b1_S7577;
      end
      test_b1_S7577: begin
        IMAGE_addr <= 7561;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S7578;
      end
      test_b1_S7578: begin
        IMAGE_addr <= 7562;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S7579;
      end
      test_b1_S7579: begin
        IMAGE_addr <= 7563;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7258;
        test_state <= test_b1_S7580;
      end
      test_b1_S7580: begin
        IMAGE_addr <= 7564;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S7581;
      end
      test_b1_S7581: begin
        IMAGE_addr <= 7565;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S7582;
      end
      test_b1_S7582: begin
        IMAGE_addr <= 7566;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7258;
        test_state <= test_b1_S7583;
      end
      test_b1_S7583: begin
        IMAGE_addr <= 7567;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S7584;
      end
      test_b1_S7584: begin
        IMAGE_addr <= 7568;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S7585;
      end
      test_b1_S7585: begin
        IMAGE_addr <= 7569;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7250;
        test_state <= test_b1_S7586;
      end
      test_b1_S7586: begin
        IMAGE_addr <= 7570;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S7587;
      end
      test_b1_S7587: begin
        IMAGE_addr <= 7571;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 16;
        test_state <= test_b1_S7588;
      end
      test_b1_S7588: begin
        IMAGE_addr <= 7572;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S7589;
      end
      test_b1_S7589: begin
        IMAGE_addr <= 7573;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7241;
        test_state <= test_b1_S7590;
      end
      test_b1_S7590: begin
        IMAGE_addr <= 7574;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S7591;
      end
      test_b1_S7591: begin
        IMAGE_addr <= 7575;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7269;
        test_state <= test_b1_S7592;
      end
      test_b1_S7592: begin
        IMAGE_addr <= 7576;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S7593;
      end
      test_b1_S7593: begin
        IMAGE_addr <= 7577;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4126;
        test_state <= test_b1_S7594;
      end
      test_b1_S7594: begin
        IMAGE_addr <= 7578;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7269;
        test_state <= test_b1_S7595;
      end
      test_b1_S7595: begin
        IMAGE_addr <= 7579;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5792;
        test_state <= test_b1_S7596;
      end
      test_b1_S7596: begin
        IMAGE_addr <= 7580;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7597;
      end
      test_b1_S7597: begin
        IMAGE_addr <= 7581;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7598;
      end
      test_b1_S7598: begin
        IMAGE_addr <= 7582;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7536;
        test_state <= test_b1_S7599;
      end
      test_b1_S7599: begin
        IMAGE_addr <= 7583;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S7600;
      end
      test_b1_S7600: begin
        IMAGE_addr <= 7584;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7594;
        test_state <= test_b1_S7601;
      end
      test_b1_S7601: begin
        IMAGE_addr <= 7585;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S7602;
      end
      test_b1_S7602: begin
        IMAGE_addr <= 7586;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S7603;
      end
      test_b1_S7603: begin
        IMAGE_addr <= 7587;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S7604;
      end
      test_b1_S7604: begin
        IMAGE_addr <= 7588;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 109;
        test_state <= test_b1_S7605;
      end
      test_b1_S7605: begin
        IMAGE_addr <= 7589;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 76;
        test_state <= test_b1_S7606;
      end
      test_b1_S7606: begin
        IMAGE_addr <= 7590;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S7607;
      end
      test_b1_S7607: begin
        IMAGE_addr <= 7591;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 102;
        test_state <= test_b1_S7608;
      end
      test_b1_S7608: begin
        IMAGE_addr <= 7592;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S7609;
      end
      test_b1_S7609: begin
        IMAGE_addr <= 7593;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7610;
      end
      test_b1_S7610: begin
        IMAGE_addr <= 7594;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7611;
      end
      test_b1_S7611: begin
        IMAGE_addr <= 7595;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7612;
      end
      test_b1_S7612: begin
        IMAGE_addr <= 7596;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S7613;
      end
      test_b1_S7613: begin
        IMAGE_addr <= 7597;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7614;
        test_state <= test_b1_S7614;
      end
      test_b1_S7614: begin
        IMAGE_addr <= 7598;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 189;
        test_state <= test_b1_S7615;
      end
      test_b1_S7615: begin
        IMAGE_addr <= 7599;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S7616;
      end
      test_b1_S7616: begin
        IMAGE_addr <= 7600;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7605;
        test_state <= test_b1_S7617;
      end
      test_b1_S7617: begin
        IMAGE_addr <= 7601;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S7618;
      end
      test_b1_S7618: begin
        IMAGE_addr <= 7602;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 32;
        test_state <= test_b1_S7619;
      end
      test_b1_S7619: begin
        IMAGE_addr <= 7603;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 790;
        test_state <= test_b1_S7620;
      end
      test_b1_S7620: begin
        IMAGE_addr <= 7604;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7621;
      end
      test_b1_S7621: begin
        IMAGE_addr <= 7605;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S7622;
      end
      test_b1_S7622: begin
        IMAGE_addr <= 7606;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7611;
        test_state <= test_b1_S7623;
      end
      test_b1_S7623: begin
        IMAGE_addr <= 7607;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S7624;
      end
      test_b1_S7624: begin
        IMAGE_addr <= 7608;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7625;
      end
      test_b1_S7625: begin
        IMAGE_addr <= 7609;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 798;
        test_state <= test_b1_S7626;
      end
      test_b1_S7626: begin
        IMAGE_addr <= 7610;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7627;
      end
      test_b1_S7627: begin
        IMAGE_addr <= 7611;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3539;
        test_state <= test_b1_S7628;
      end
      test_b1_S7628: begin
        IMAGE_addr <= 7612;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 20;
        test_state <= test_b1_S7629;
      end
      test_b1_S7629: begin
        IMAGE_addr <= 7613;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7630;
      end
      test_b1_S7630: begin
        IMAGE_addr <= 7614;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3433;
        test_state <= test_b1_S7631;
      end
      test_b1_S7631: begin
        IMAGE_addr <= 7615;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 27;
        test_state <= test_b1_S7632;
      end
      test_b1_S7632: begin
        IMAGE_addr <= 7616;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7633;
      end
      test_b1_S7633: begin
        IMAGE_addr <= 7617;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7634;
      end
      test_b1_S7634: begin
        IMAGE_addr <= 7618;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7582;
        test_state <= test_b1_S7635;
      end
      test_b1_S7635: begin
        IMAGE_addr <= 7619;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S7636;
      end
      test_b1_S7636: begin
        IMAGE_addr <= 7620;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7631;
        test_state <= test_b1_S7637;
      end
      test_b1_S7637: begin
        IMAGE_addr <= 7621;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S7638;
      end
      test_b1_S7638: begin
        IMAGE_addr <= 7622;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S7639;
      end
      test_b1_S7639: begin
        IMAGE_addr <= 7623;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S7640;
      end
      test_b1_S7640: begin
        IMAGE_addr <= 7624;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 109;
        test_state <= test_b1_S7641;
      end
      test_b1_S7641: begin
        IMAGE_addr <= 7625;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 82;
        test_state <= test_b1_S7642;
      end
      test_b1_S7642: begin
        IMAGE_addr <= 7626;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S7643;
      end
      test_b1_S7643: begin
        IMAGE_addr <= 7627;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 103;
        test_state <= test_b1_S7644;
      end
      test_b1_S7644: begin
        IMAGE_addr <= 7628;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 104;
        test_state <= test_b1_S7645;
      end
      test_b1_S7645: begin
        IMAGE_addr <= 7629;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S7646;
      end
      test_b1_S7646: begin
        IMAGE_addr <= 7630;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7647;
      end
      test_b1_S7647: begin
        IMAGE_addr <= 7631;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7648;
      end
      test_b1_S7648: begin
        IMAGE_addr <= 7632;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7649;
      end
      test_b1_S7649: begin
        IMAGE_addr <= 7633;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7269;
        test_state <= test_b1_S7650;
      end
      test_b1_S7650: begin
        IMAGE_addr <= 7634;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S7651;
      end
      test_b1_S7651: begin
        IMAGE_addr <= 7635;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7641;
        test_state <= test_b1_S7652;
      end
      test_b1_S7652: begin
        IMAGE_addr <= 7636;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S7653;
      end
      test_b1_S7653: begin
        IMAGE_addr <= 7637;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7654;
      end
      test_b1_S7654: begin
        IMAGE_addr <= 7638;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 909;
        test_state <= test_b1_S7655;
      end
      test_b1_S7655: begin
        IMAGE_addr <= 7639;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4148;
        test_state <= test_b1_S7656;
      end
      test_b1_S7656: begin
        IMAGE_addr <= 7640;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7657;
      end
      test_b1_S7657: begin
        IMAGE_addr <= 7641;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S7658;
      end
      test_b1_S7658: begin
        IMAGE_addr <= 7642;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7647;
        test_state <= test_b1_S7659;
      end
      test_b1_S7659: begin
        IMAGE_addr <= 7643;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 132;
        test_state <= test_b1_S7660;
      end
      test_b1_S7660: begin
        IMAGE_addr <= 7644;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 877;
        test_state <= test_b1_S7661;
      end
      test_b1_S7661: begin
        IMAGE_addr <= 7645;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4126;
        test_state <= test_b1_S7662;
      end
      test_b1_S7662: begin
        IMAGE_addr <= 7646;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7663;
      end
      test_b1_S7663: begin
        IMAGE_addr <= 7647;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S7664;
      end
      test_b1_S7664: begin
        IMAGE_addr <= 7648;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7651;
        test_state <= test_b1_S7665;
      end
      test_b1_S7665: begin
        IMAGE_addr <= 7649;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7289;
        test_state <= test_b1_S7666;
      end
      test_b1_S7666: begin
        IMAGE_addr <= 7650;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7667;
      end
      test_b1_S7667: begin
        IMAGE_addr <= 7651;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3582;
        test_state <= test_b1_S7668;
      end
      test_b1_S7668: begin
        IMAGE_addr <= 7652;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5792;
        test_state <= test_b1_S7669;
      end
      test_b1_S7669: begin
        IMAGE_addr <= 7653;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7670;
      end
      test_b1_S7670: begin
        IMAGE_addr <= 7654;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7671;
      end
      test_b1_S7671: begin
        IMAGE_addr <= 7655;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7618;
        test_state <= test_b1_S7672;
      end
      test_b1_S7672: begin
        IMAGE_addr <= 7656;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S7673;
      end
      test_b1_S7673: begin
        IMAGE_addr <= 7657;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7666;
        test_state <= test_b1_S7674;
      end
      test_b1_S7674: begin
        IMAGE_addr <= 7658;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 112;
        test_state <= test_b1_S7675;
      end
      test_b1_S7675: begin
        IMAGE_addr <= 7659;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S7676;
      end
      test_b1_S7676: begin
        IMAGE_addr <= 7660;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S7677;
      end
      test_b1_S7677: begin
        IMAGE_addr <= 7661;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 112;
        test_state <= test_b1_S7678;
      end
      test_b1_S7678: begin
        IMAGE_addr <= 7662;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S7679;
      end
      test_b1_S7679: begin
        IMAGE_addr <= 7663;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 110;
        test_state <= test_b1_S7680;
      end
      test_b1_S7680: begin
        IMAGE_addr <= 7664;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 100;
        test_state <= test_b1_S7681;
      end
      test_b1_S7681: begin
        IMAGE_addr <= 7665;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7682;
      end
      test_b1_S7682: begin
        IMAGE_addr <= 7666;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7683;
      end
      test_b1_S7683: begin
        IMAGE_addr <= 7667;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7684;
      end
      test_b1_S7684: begin
        IMAGE_addr <= 7668;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7269;
        test_state <= test_b1_S7685;
      end
      test_b1_S7685: begin
        IMAGE_addr <= 7669;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S7686;
      end
      test_b1_S7686: begin
        IMAGE_addr <= 7670;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7687;
      end
      test_b1_S7687: begin
        IMAGE_addr <= 7671;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 909;
        test_state <= test_b1_S7688;
      end
      test_b1_S7688: begin
        IMAGE_addr <= 7672;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4148;
        test_state <= test_b1_S7689;
      end
      test_b1_S7689: begin
        IMAGE_addr <= 7673;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 886;
        test_state <= test_b1_S7690;
      end
      test_b1_S7690: begin
        IMAGE_addr <= 7674;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7269;
        test_state <= test_b1_S7691;
      end
      test_b1_S7691: begin
        IMAGE_addr <= 7675;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S7692;
      end
      test_b1_S7692: begin
        IMAGE_addr <= 7676;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S7693;
      end
      test_b1_S7693: begin
        IMAGE_addr <= 7677;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4126;
        test_state <= test_b1_S7694;
      end
      test_b1_S7694: begin
        IMAGE_addr <= 7678;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 774;
        test_state <= test_b1_S7695;
      end
      test_b1_S7695: begin
        IMAGE_addr <= 7679;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S7696;
      end
      test_b1_S7696: begin
        IMAGE_addr <= 7680;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 886;
        test_state <= test_b1_S7697;
      end
      test_b1_S7697: begin
        IMAGE_addr <= 7681;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 766;
        test_state <= test_b1_S7698;
      end
      test_b1_S7698: begin
        IMAGE_addr <= 7682;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7269;
        test_state <= test_b1_S7699;
      end
      test_b1_S7699: begin
        IMAGE_addr <= 7683;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 16;
        test_state <= test_b1_S7700;
      end
      test_b1_S7700: begin
        IMAGE_addr <= 7684;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S7701;
      end
      test_b1_S7701: begin
        IMAGE_addr <= 7685;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4126;
        test_state <= test_b1_S7702;
      end
      test_b1_S7702: begin
        IMAGE_addr <= 7686;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7269;
        test_state <= test_b1_S7703;
      end
      test_b1_S7703: begin
        IMAGE_addr <= 7687;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5792;
        test_state <= test_b1_S7704;
      end
      test_b1_S7704: begin
        IMAGE_addr <= 7688;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7705;
      end
      test_b1_S7705: begin
        IMAGE_addr <= 7689;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7706;
      end
      test_b1_S7706: begin
        IMAGE_addr <= 7690;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7655;
        test_state <= test_b1_S7707;
      end
      test_b1_S7707: begin
        IMAGE_addr <= 7691;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S7708;
      end
      test_b1_S7708: begin
        IMAGE_addr <= 7692;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7700;
        test_state <= test_b1_S7709;
      end
      test_b1_S7709: begin
        IMAGE_addr <= 7693;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S7710;
      end
      test_b1_S7710: begin
        IMAGE_addr <= 7694;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 112;
        test_state <= test_b1_S7711;
      end
      test_b1_S7711: begin
        IMAGE_addr <= 7695;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 112;
        test_state <= test_b1_S7712;
      end
      test_b1_S7712: begin
        IMAGE_addr <= 7696;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S7713;
      end
      test_b1_S7713: begin
        IMAGE_addr <= 7697;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 110;
        test_state <= test_b1_S7714;
      end
      test_b1_S7714: begin
        IMAGE_addr <= 7698;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 100;
        test_state <= test_b1_S7715;
      end
      test_b1_S7715: begin
        IMAGE_addr <= 7699;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7716;
      end
      test_b1_S7716: begin
        IMAGE_addr <= 7700;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7717;
      end
      test_b1_S7717: begin
        IMAGE_addr <= 7701;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7718;
      end
      test_b1_S7718: begin
        IMAGE_addr <= 7702;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S7719;
      end
      test_b1_S7719: begin
        IMAGE_addr <= 7703;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7666;
        test_state <= test_b1_S7720;
      end
      test_b1_S7720: begin
        IMAGE_addr <= 7704;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7721;
      end
      test_b1_S7721: begin
        IMAGE_addr <= 7705;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7722;
      end
      test_b1_S7722: begin
        IMAGE_addr <= 7706;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7690;
        test_state <= test_b1_S7723;
      end
      test_b1_S7723: begin
        IMAGE_addr <= 7707;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S7724;
      end
      test_b1_S7724: begin
        IMAGE_addr <= 7708;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7720;
        test_state <= test_b1_S7725;
      end
      test_b1_S7725: begin
        IMAGE_addr <= 7709;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S7726;
      end
      test_b1_S7726: begin
        IMAGE_addr <= 7710;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 112;
        test_state <= test_b1_S7727;
      end
      test_b1_S7727: begin
        IMAGE_addr <= 7711;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 112;
        test_state <= test_b1_S7728;
      end
      test_b1_S7728: begin
        IMAGE_addr <= 7712;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S7729;
      end
      test_b1_S7729: begin
        IMAGE_addr <= 7713;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 110;
        test_state <= test_b1_S7730;
      end
      test_b1_S7730: begin
        IMAGE_addr <= 7714;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 100;
        test_state <= test_b1_S7731;
      end
      test_b1_S7731: begin
        IMAGE_addr <= 7715;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 67;
        test_state <= test_b1_S7732;
      end
      test_b1_S7732: begin
        IMAGE_addr <= 7716;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 104;
        test_state <= test_b1_S7733;
      end
      test_b1_S7733: begin
        IMAGE_addr <= 7717;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S7734;
      end
      test_b1_S7734: begin
        IMAGE_addr <= 7718;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S7735;
      end
      test_b1_S7735: begin
        IMAGE_addr <= 7719;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7736;
      end
      test_b1_S7736: begin
        IMAGE_addr <= 7720;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7737;
      end
      test_b1_S7737: begin
        IMAGE_addr <= 7721;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7738;
      end
      test_b1_S7738: begin
        IMAGE_addr <= 7722;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S7739;
      end
      test_b1_S7739: begin
        IMAGE_addr <= 7723;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5792;
        test_state <= test_b1_S7740;
      end
      test_b1_S7740: begin
        IMAGE_addr <= 7724;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S7741;
      end
      test_b1_S7741: begin
        IMAGE_addr <= 7725;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7734;
        test_state <= test_b1_S7742;
      end
      test_b1_S7742: begin
        IMAGE_addr <= 7726;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 886;
        test_state <= test_b1_S7743;
      end
      test_b1_S7743: begin
        IMAGE_addr <= 7727;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 16;
        test_state <= test_b1_S7744;
      end
      test_b1_S7744: begin
        IMAGE_addr <= 7728;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 197;
        test_state <= test_b1_S7745;
      end
      test_b1_S7745: begin
        IMAGE_addr <= 7729;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S7746;
      end
      test_b1_S7746: begin
        IMAGE_addr <= 7730;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7747;
      end
      test_b1_S7747: begin
        IMAGE_addr <= 7731;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S7748;
      end
      test_b1_S7748: begin
        IMAGE_addr <= 7732;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S7749;
      end
      test_b1_S7749: begin
        IMAGE_addr <= 7733;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7750;
      end
      test_b1_S7750: begin
        IMAGE_addr <= 7734;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 774;
        test_state <= test_b1_S7751;
      end
      test_b1_S7751: begin
        IMAGE_addr <= 7735;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7752;
      end
      test_b1_S7752: begin
        IMAGE_addr <= 7736;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7753;
      end
      test_b1_S7753: begin
        IMAGE_addr <= 7737;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7706;
        test_state <= test_b1_S7754;
      end
      test_b1_S7754: begin
        IMAGE_addr <= 7738;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S7755;
      end
      test_b1_S7755: begin
        IMAGE_addr <= 7739;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7748;
        test_state <= test_b1_S7756;
      end
      test_b1_S7756: begin
        IMAGE_addr <= 7740;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S7757;
      end
      test_b1_S7757: begin
        IMAGE_addr <= 7741;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 111;
        test_state <= test_b1_S7758;
      end
      test_b1_S7758: begin
        IMAGE_addr <= 7742;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 76;
        test_state <= test_b1_S7759;
      end
      test_b1_S7759: begin
        IMAGE_addr <= 7743;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 111;
        test_state <= test_b1_S7760;
      end
      test_b1_S7760: begin
        IMAGE_addr <= 7744;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 119;
        test_state <= test_b1_S7761;
      end
      test_b1_S7761: begin
        IMAGE_addr <= 7745;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S7762;
      end
      test_b1_S7762: begin
        IMAGE_addr <= 7746;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S7763;
      end
      test_b1_S7763: begin
        IMAGE_addr <= 7747;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7764;
      end
      test_b1_S7764: begin
        IMAGE_addr <= 7748;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7765;
      end
      test_b1_S7765: begin
        IMAGE_addr <= 7749;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7766;
      end
      test_b1_S7766: begin
        IMAGE_addr <= 7750;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 886;
        test_state <= test_b1_S7767;
      end
      test_b1_S7767: begin
        IMAGE_addr <= 7751;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 26;
        test_state <= test_b1_S7768;
      end
      test_b1_S7768: begin
        IMAGE_addr <= 7752;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S7769;
      end
      test_b1_S7769: begin
        IMAGE_addr <= 7753;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7779;
        test_state <= test_b1_S7770;
      end
      test_b1_S7770: begin
        IMAGE_addr <= 7754;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7269;
        test_state <= test_b1_S7771;
      end
      test_b1_S7771: begin
        IMAGE_addr <= 7755;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 16;
        test_state <= test_b1_S7772;
      end
      test_b1_S7772: begin
        IMAGE_addr <= 7756;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S7773;
      end
      test_b1_S7773: begin
        IMAGE_addr <= 7757;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7776;
        test_state <= test_b1_S7774;
      end
      test_b1_S7774: begin
        IMAGE_addr <= 7758;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 189;
        test_state <= test_b1_S7775;
      end
      test_b1_S7775: begin
        IMAGE_addr <= 7759;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S7776;
      end
      test_b1_S7776: begin
        IMAGE_addr <= 7760;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S7777;
      end
      test_b1_S7777: begin
        IMAGE_addr <= 7761;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 65;
        test_state <= test_b1_S7778;
      end
      test_b1_S7778: begin
        IMAGE_addr <= 7762;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S7779;
      end
      test_b1_S7779: begin
        IMAGE_addr <= 7763;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 90;
        test_state <= test_b1_S7780;
      end
      test_b1_S7780: begin
        IMAGE_addr <= 7764;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4214;
        test_state <= test_b1_S7781;
      end
      test_b1_S7781: begin
        IMAGE_addr <= 7765;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S7782;
      end
      test_b1_S7782: begin
        IMAGE_addr <= 7766;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7774;
        test_state <= test_b1_S7783;
      end
      test_b1_S7783: begin
        IMAGE_addr <= 7767;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S7784;
      end
      test_b1_S7784: begin
        IMAGE_addr <= 7768;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S7785;
      end
      test_b1_S7785: begin
        IMAGE_addr <= 7769;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 16;
        test_state <= test_b1_S7786;
      end
      test_b1_S7786: begin
        IMAGE_addr <= 7770;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S7787;
      end
      test_b1_S7787: begin
        IMAGE_addr <= 7771;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 65;
        test_state <= test_b1_S7788;
      end
      test_b1_S7788: begin
        IMAGE_addr <= 7772;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 17;
        test_state <= test_b1_S7789;
      end
      test_b1_S7789: begin
        IMAGE_addr <= 7773;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7790;
      end
      test_b1_S7790: begin
        IMAGE_addr <= 7774;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 751;
        test_state <= test_b1_S7791;
      end
      test_b1_S7791: begin
        IMAGE_addr <= 7775;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7792;
      end
      test_b1_S7792: begin
        IMAGE_addr <= 7776;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 766;
        test_state <= test_b1_S7793;
      end
      test_b1_S7793: begin
        IMAGE_addr <= 7777;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S7794;
      end
      test_b1_S7794: begin
        IMAGE_addr <= 7778;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7795;
      end
      test_b1_S7795: begin
        IMAGE_addr <= 7779;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3912;
        test_state <= test_b1_S7796;
      end
      test_b1_S7796: begin
        IMAGE_addr <= 7780;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S7797;
      end
      test_b1_S7797: begin
        IMAGE_addr <= 7781;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7269;
        test_state <= test_b1_S7798;
      end
      test_b1_S7798: begin
        IMAGE_addr <= 7782;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5792;
        test_state <= test_b1_S7799;
      end
      test_b1_S7799: begin
        IMAGE_addr <= 7783;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7800;
      end
      test_b1_S7800: begin
        IMAGE_addr <= 7784;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7801;
      end
      test_b1_S7801: begin
        IMAGE_addr <= 7785;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7737;
        test_state <= test_b1_S7802;
      end
      test_b1_S7802: begin
        IMAGE_addr <= 7786;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S7803;
      end
      test_b1_S7803: begin
        IMAGE_addr <= 7787;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7796;
        test_state <= test_b1_S7804;
      end
      test_b1_S7804: begin
        IMAGE_addr <= 7788;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S7805;
      end
      test_b1_S7805: begin
        IMAGE_addr <= 7789;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 111;
        test_state <= test_b1_S7806;
      end
      test_b1_S7806: begin
        IMAGE_addr <= 7790;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 85;
        test_state <= test_b1_S7807;
      end
      test_b1_S7807: begin
        IMAGE_addr <= 7791;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 112;
        test_state <= test_b1_S7808;
      end
      test_b1_S7808: begin
        IMAGE_addr <= 7792;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 112;
        test_state <= test_b1_S7809;
      end
      test_b1_S7809: begin
        IMAGE_addr <= 7793;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S7810;
      end
      test_b1_S7810: begin
        IMAGE_addr <= 7794;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S7811;
      end
      test_b1_S7811: begin
        IMAGE_addr <= 7795;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7812;
      end
      test_b1_S7812: begin
        IMAGE_addr <= 7796;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7813;
      end
      test_b1_S7813: begin
        IMAGE_addr <= 7797;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7814;
      end
      test_b1_S7814: begin
        IMAGE_addr <= 7798;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 886;
        test_state <= test_b1_S7815;
      end
      test_b1_S7815: begin
        IMAGE_addr <= 7799;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 26;
        test_state <= test_b1_S7816;
      end
      test_b1_S7816: begin
        IMAGE_addr <= 7800;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S7817;
      end
      test_b1_S7817: begin
        IMAGE_addr <= 7801;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7827;
        test_state <= test_b1_S7818;
      end
      test_b1_S7818: begin
        IMAGE_addr <= 7802;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7269;
        test_state <= test_b1_S7819;
      end
      test_b1_S7819: begin
        IMAGE_addr <= 7803;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 16;
        test_state <= test_b1_S7820;
      end
      test_b1_S7820: begin
        IMAGE_addr <= 7804;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S7821;
      end
      test_b1_S7821: begin
        IMAGE_addr <= 7805;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7824;
        test_state <= test_b1_S7822;
      end
      test_b1_S7822: begin
        IMAGE_addr <= 7806;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 189;
        test_state <= test_b1_S7823;
      end
      test_b1_S7823: begin
        IMAGE_addr <= 7807;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S7824;
      end
      test_b1_S7824: begin
        IMAGE_addr <= 7808;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S7825;
      end
      test_b1_S7825: begin
        IMAGE_addr <= 7809;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S7826;
      end
      test_b1_S7826: begin
        IMAGE_addr <= 7810;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S7827;
      end
      test_b1_S7827: begin
        IMAGE_addr <= 7811;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 122;
        test_state <= test_b1_S7828;
      end
      test_b1_S7828: begin
        IMAGE_addr <= 7812;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4214;
        test_state <= test_b1_S7829;
      end
      test_b1_S7829: begin
        IMAGE_addr <= 7813;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S7830;
      end
      test_b1_S7830: begin
        IMAGE_addr <= 7814;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7822;
        test_state <= test_b1_S7831;
      end
      test_b1_S7831: begin
        IMAGE_addr <= 7815;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S7832;
      end
      test_b1_S7832: begin
        IMAGE_addr <= 7816;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 65;
        test_state <= test_b1_S7833;
      end
      test_b1_S7833: begin
        IMAGE_addr <= 7817;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 16;
        test_state <= test_b1_S7834;
      end
      test_b1_S7834: begin
        IMAGE_addr <= 7818;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S7835;
      end
      test_b1_S7835: begin
        IMAGE_addr <= 7819;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S7836;
      end
      test_b1_S7836: begin
        IMAGE_addr <= 7820;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 17;
        test_state <= test_b1_S7837;
      end
      test_b1_S7837: begin
        IMAGE_addr <= 7821;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7838;
      end
      test_b1_S7838: begin
        IMAGE_addr <= 7822;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 751;
        test_state <= test_b1_S7839;
      end
      test_b1_S7839: begin
        IMAGE_addr <= 7823;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7840;
      end
      test_b1_S7840: begin
        IMAGE_addr <= 7824;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 766;
        test_state <= test_b1_S7841;
      end
      test_b1_S7841: begin
        IMAGE_addr <= 7825;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S7842;
      end
      test_b1_S7842: begin
        IMAGE_addr <= 7826;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7843;
      end
      test_b1_S7843: begin
        IMAGE_addr <= 7827;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3912;
        test_state <= test_b1_S7844;
      end
      test_b1_S7844: begin
        IMAGE_addr <= 7828;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S7845;
      end
      test_b1_S7845: begin
        IMAGE_addr <= 7829;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7269;
        test_state <= test_b1_S7846;
      end
      test_b1_S7846: begin
        IMAGE_addr <= 7830;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5792;
        test_state <= test_b1_S7847;
      end
      test_b1_S7847: begin
        IMAGE_addr <= 7831;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7848;
      end
      test_b1_S7848: begin
        IMAGE_addr <= 7832;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7849;
      end
      test_b1_S7849: begin
        IMAGE_addr <= 7833;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7785;
        test_state <= test_b1_S7850;
      end
      test_b1_S7850: begin
        IMAGE_addr <= 7834;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S7851;
      end
      test_b1_S7851: begin
        IMAGE_addr <= 7835;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7844;
        test_state <= test_b1_S7852;
      end
      test_b1_S7852: begin
        IMAGE_addr <= 7836;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S7853;
      end
      test_b1_S7853: begin
        IMAGE_addr <= 7837;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S7854;
      end
      test_b1_S7854: begin
        IMAGE_addr <= 7838;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 118;
        test_state <= test_b1_S7855;
      end
      test_b1_S7855: begin
        IMAGE_addr <= 7839;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S7856;
      end
      test_b1_S7856: begin
        IMAGE_addr <= 7840;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S7857;
      end
      test_b1_S7857: begin
        IMAGE_addr <= 7841;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S7858;
      end
      test_b1_S7858: begin
        IMAGE_addr <= 7842;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S7859;
      end
      test_b1_S7859: begin
        IMAGE_addr <= 7843;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7860;
      end
      test_b1_S7860: begin
        IMAGE_addr <= 7844;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7861;
      end
      test_b1_S7861: begin
        IMAGE_addr <= 7845;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7862;
      end
      test_b1_S7862: begin
        IMAGE_addr <= 7846;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S7863;
      end
      test_b1_S7863: begin
        IMAGE_addr <= 7847;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5792;
        test_state <= test_b1_S7864;
      end
      test_b1_S7864: begin
        IMAGE_addr <= 7848;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7164;
        test_state <= test_b1_S7865;
      end
      test_b1_S7865: begin
        IMAGE_addr <= 7849;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S7866;
      end
      test_b1_S7866: begin
        IMAGE_addr <= 7850;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 877;
        test_state <= test_b1_S7867;
      end
      test_b1_S7867: begin
        IMAGE_addr <= 7851;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S7868;
      end
      test_b1_S7868: begin
        IMAGE_addr <= 7852;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7857;
        test_state <= test_b1_S7869;
      end
      test_b1_S7869: begin
        IMAGE_addr <= 7853;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 886;
        test_state <= test_b1_S7870;
      end
      test_b1_S7870: begin
        IMAGE_addr <= 7854;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 16;
        test_state <= test_b1_S7871;
      end
      test_b1_S7871: begin
        IMAGE_addr <= 7855;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 27;
        test_state <= test_b1_S7872;
      end
      test_b1_S7872: begin
        IMAGE_addr <= 7856;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7873;
      end
      test_b1_S7873: begin
        IMAGE_addr <= 7857;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3539;
        test_state <= test_b1_S7874;
      end
      test_b1_S7874: begin
        IMAGE_addr <= 7858;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S7875;
      end
      test_b1_S7875: begin
        IMAGE_addr <= 7859;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S7876;
      end
      test_b1_S7876: begin
        IMAGE_addr <= 7860;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7866;
        test_state <= test_b1_S7877;
      end
      test_b1_S7877: begin
        IMAGE_addr <= 7861;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S7878;
      end
      test_b1_S7878: begin
        IMAGE_addr <= 7862;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S7879;
      end
      test_b1_S7879: begin
        IMAGE_addr <= 7863;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7097;
        test_state <= test_b1_S7880;
      end
      test_b1_S7880: begin
        IMAGE_addr <= 7864;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 27;
        test_state <= test_b1_S7881;
      end
      test_b1_S7881: begin
        IMAGE_addr <= 7865;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7882;
      end
      test_b1_S7882: begin
        IMAGE_addr <= 7866;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3841;
        test_state <= test_b1_S7883;
      end
      test_b1_S7883: begin
        IMAGE_addr <= 7867;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S7884;
      end
      test_b1_S7884: begin
        IMAGE_addr <= 7868;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7069;
        test_state <= test_b1_S7885;
      end
      test_b1_S7885: begin
        IMAGE_addr <= 7869;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5792;
        test_state <= test_b1_S7886;
      end
      test_b1_S7886: begin
        IMAGE_addr <= 7870;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7887;
      end
      test_b1_S7887: begin
        IMAGE_addr <= 7871;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7888;
      end
      test_b1_S7888: begin
        IMAGE_addr <= 7872;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7833;
        test_state <= test_b1_S7889;
      end
      test_b1_S7889: begin
        IMAGE_addr <= 7873;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S7890;
      end
      test_b1_S7890: begin
        IMAGE_addr <= 7874;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7881;
        test_state <= test_b1_S7891;
      end
      test_b1_S7891: begin
        IMAGE_addr <= 7875;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S7892;
      end
      test_b1_S7892: begin
        IMAGE_addr <= 7876;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 112;
        test_state <= test_b1_S7893;
      end
      test_b1_S7893: begin
        IMAGE_addr <= 7877;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 108;
        test_state <= test_b1_S7894;
      end
      test_b1_S7894: begin
        IMAGE_addr <= 7878;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S7895;
      end
      test_b1_S7895: begin
        IMAGE_addr <= 7879;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S7896;
      end
      test_b1_S7896: begin
        IMAGE_addr <= 7880;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7897;
      end
      test_b1_S7897: begin
        IMAGE_addr <= 7881;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7898;
      end
      test_b1_S7898: begin
        IMAGE_addr <= 7882;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7899;
      end
      test_b1_S7899: begin
        IMAGE_addr <= 7883;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 132;
        test_state <= test_b1_S7900;
      end
      test_b1_S7900: begin
        IMAGE_addr <= 7884;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 132;
        test_state <= test_b1_S7901;
      end
      test_b1_S7901: begin
        IMAGE_addr <= 7885;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S7902;
      end
      test_b1_S7902: begin
        IMAGE_addr <= 7886;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7903;
      end
      test_b1_S7903: begin
        IMAGE_addr <= 7887;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S7904;
      end
      test_b1_S7904: begin
        IMAGE_addr <= 7888;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7549;
        test_state <= test_b1_S7905;
      end
      test_b1_S7905: begin
        IMAGE_addr <= 7889;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S7906;
      end
      test_b1_S7906: begin
        IMAGE_addr <= 7890;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7893;
        test_state <= test_b1_S7907;
      end
      test_b1_S7907: begin
        IMAGE_addr <= 7891;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 16;
        test_state <= test_b1_S7908;
      end
      test_b1_S7908: begin
        IMAGE_addr <= 7892;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7909;
      end
      test_b1_S7909: begin
        IMAGE_addr <= 7893;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 766;
        test_state <= test_b1_S7910;
      end
      test_b1_S7910: begin
        IMAGE_addr <= 7894;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7911;
      end
      test_b1_S7911: begin
        IMAGE_addr <= 7895;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7912;
      end
      test_b1_S7912: begin
        IMAGE_addr <= 7896;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7872;
        test_state <= test_b1_S7913;
      end
      test_b1_S7913: begin
        IMAGE_addr <= 7897;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S7914;
      end
      test_b1_S7914: begin
        IMAGE_addr <= 7898;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7911;
        test_state <= test_b1_S7915;
      end
      test_b1_S7915: begin
        IMAGE_addr <= 7899;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S7916;
      end
      test_b1_S7916: begin
        IMAGE_addr <= 7900;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 112;
        test_state <= test_b1_S7917;
      end
      test_b1_S7917: begin
        IMAGE_addr <= 7901;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 108;
        test_state <= test_b1_S7918;
      end
      test_b1_S7918: begin
        IMAGE_addr <= 7902;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S7919;
      end
      test_b1_S7919: begin
        IMAGE_addr <= 7903;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S7920;
      end
      test_b1_S7920: begin
        IMAGE_addr <= 7904;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 65;
        test_state <= test_b1_S7921;
      end
      test_b1_S7921: begin
        IMAGE_addr <= 7905;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S7922;
      end
      test_b1_S7922: begin
        IMAGE_addr <= 7906;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 67;
        test_state <= test_b1_S7923;
      end
      test_b1_S7923: begin
        IMAGE_addr <= 7907;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 104;
        test_state <= test_b1_S7924;
      end
      test_b1_S7924: begin
        IMAGE_addr <= 7908;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S7925;
      end
      test_b1_S7925: begin
        IMAGE_addr <= 7909;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S7926;
      end
      test_b1_S7926: begin
        IMAGE_addr <= 7910;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7927;
      end
      test_b1_S7927: begin
        IMAGE_addr <= 7911;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7928;
      end
      test_b1_S7928: begin
        IMAGE_addr <= 7912;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7929;
      end
      test_b1_S7929: begin
        IMAGE_addr <= 7913;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 132;
        test_state <= test_b1_S7930;
      end
      test_b1_S7930: begin
        IMAGE_addr <= 7914;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 132;
        test_state <= test_b1_S7931;
      end
      test_b1_S7931: begin
        IMAGE_addr <= 7915;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 132;
        test_state <= test_b1_S7932;
      end
      test_b1_S7932: begin
        IMAGE_addr <= 7916;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S7933;
      end
      test_b1_S7933: begin
        IMAGE_addr <= 7917;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7466;
        test_state <= test_b1_S7934;
      end
      test_b1_S7934: begin
        IMAGE_addr <= 7918;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 132;
        test_state <= test_b1_S7935;
      end
      test_b1_S7935: begin
        IMAGE_addr <= 7919;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 17;
        test_state <= test_b1_S7936;
      end
      test_b1_S7936: begin
        IMAGE_addr <= 7920;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 26;
        test_state <= test_b1_S7937;
      end
      test_b1_S7937: begin
        IMAGE_addr <= 7921;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S7938;
      end
      test_b1_S7938: begin
        IMAGE_addr <= 7922;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7939;
      end
      test_b1_S7939: begin
        IMAGE_addr <= 7923;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S7940;
      end
      test_b1_S7940: begin
        IMAGE_addr <= 7924;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7549;
        test_state <= test_b1_S7941;
      end
      test_b1_S7941: begin
        IMAGE_addr <= 7925;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S7942;
      end
      test_b1_S7942: begin
        IMAGE_addr <= 7926;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7930;
        test_state <= test_b1_S7943;
      end
      test_b1_S7943: begin
        IMAGE_addr <= 7927;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7466;
        test_state <= test_b1_S7944;
      end
      test_b1_S7944: begin
        IMAGE_addr <= 7928;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 26;
        test_state <= test_b1_S7945;
      end
      test_b1_S7945: begin
        IMAGE_addr <= 7929;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7946;
      end
      test_b1_S7946: begin
        IMAGE_addr <= 7930;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 766;
        test_state <= test_b1_S7947;
      end
      test_b1_S7947: begin
        IMAGE_addr <= 7931;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7948;
      end
      test_b1_S7948: begin
        IMAGE_addr <= 7932;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7949;
      end
      test_b1_S7949: begin
        IMAGE_addr <= 7933;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7896;
        test_state <= test_b1_S7950;
      end
      test_b1_S7950: begin
        IMAGE_addr <= 7934;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 306;
        test_state <= test_b1_S7951;
      end
      test_b1_S7951: begin
        IMAGE_addr <= 7935;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7949;
        test_state <= test_b1_S7952;
      end
      test_b1_S7952: begin
        IMAGE_addr <= 7936;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S7953;
      end
      test_b1_S7953: begin
        IMAGE_addr <= 7937;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 112;
        test_state <= test_b1_S7954;
      end
      test_b1_S7954: begin
        IMAGE_addr <= 7938;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 108;
        test_state <= test_b1_S7955;
      end
      test_b1_S7955: begin
        IMAGE_addr <= 7939;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S7956;
      end
      test_b1_S7956: begin
        IMAGE_addr <= 7940;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S7957;
      end
      test_b1_S7957: begin
        IMAGE_addr <= 7941;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 65;
        test_state <= test_b1_S7958;
      end
      test_b1_S7958: begin
        IMAGE_addr <= 7942;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S7959;
      end
      test_b1_S7959: begin
        IMAGE_addr <= 7943;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 67;
        test_state <= test_b1_S7960;
      end
      test_b1_S7960: begin
        IMAGE_addr <= 7944;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 104;
        test_state <= test_b1_S7961;
      end
      test_b1_S7961: begin
        IMAGE_addr <= 7945;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S7962;
      end
      test_b1_S7962: begin
        IMAGE_addr <= 7946;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S7963;
      end
      test_b1_S7963: begin
        IMAGE_addr <= 7947;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 58;
        test_state <= test_b1_S7964;
      end
      test_b1_S7964: begin
        IMAGE_addr <= 7948;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7965;
      end
      test_b1_S7965: begin
        IMAGE_addr <= 7949;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7966;
      end
      test_b1_S7966: begin
        IMAGE_addr <= 7950;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7967;
      end
      test_b1_S7967: begin
        IMAGE_addr <= 7951;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S7968;
      end
      test_b1_S7968: begin
        IMAGE_addr <= 7952;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 32;
        test_state <= test_b1_S7969;
      end
      test_b1_S7969: begin
        IMAGE_addr <= 7953;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 562;
        test_state <= test_b1_S7970;
      end
      test_b1_S7970: begin
        IMAGE_addr <= 7954;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 400;
        test_state <= test_b1_S7971;
      end
      test_b1_S7971: begin
        IMAGE_addr <= 7955;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S7972;
      end
      test_b1_S7972: begin
        IMAGE_addr <= 7956;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 310;
        test_state <= test_b1_S7973;
      end
      test_b1_S7973: begin
        IMAGE_addr <= 7957;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S7974;
      end
      test_b1_S7974: begin
        IMAGE_addr <= 7958;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7911;
        test_state <= test_b1_S7975;
      end
      test_b1_S7975: begin
        IMAGE_addr <= 7959;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S7976;
      end
      test_b1_S7976: begin
        IMAGE_addr <= 7960;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7977;
      end
      test_b1_S7977: begin
        IMAGE_addr <= 7961;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S7978;
      end
      test_b1_S7978: begin
        IMAGE_addr <= 7962;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7172;
        test_state <= test_b1_S7979;
      end
      test_b1_S7979: begin
        IMAGE_addr <= 7963;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4705;
        test_state <= test_b1_S7980;
      end
      test_b1_S7980: begin
        IMAGE_addr <= 7964;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7969;
        test_state <= test_b1_S7981;
      end
      test_b1_S7981: begin
        IMAGE_addr <= 7965;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 95;
        test_state <= test_b1_S7982;
      end
      test_b1_S7982: begin
        IMAGE_addr <= 7966;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 95;
        test_state <= test_b1_S7983;
      end
      test_b1_S7983: begin
        IMAGE_addr <= 7967;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 94;
        test_state <= test_b1_S7984;
      end
      test_b1_S7984: begin
        IMAGE_addr <= 7968;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7985;
      end
      test_b1_S7985: begin
        IMAGE_addr <= 7969;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7986;
      end
      test_b1_S7986: begin
        IMAGE_addr <= 7970;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S7987;
      end
      test_b1_S7987: begin
        IMAGE_addr <= 7971;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S7988;
      end
      test_b1_S7988: begin
        IMAGE_addr <= 7972;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 39;
        test_state <= test_b1_S7989;
      end
      test_b1_S7989: begin
        IMAGE_addr <= 7973;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7911;
        test_state <= test_b1_S7990;
      end
      test_b1_S7990: begin
        IMAGE_addr <= 7974;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1232;
        test_state <= test_b1_S7991;
      end
      test_b1_S7991: begin
        IMAGE_addr <= 7975;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S7992;
      end
      test_b1_S7992: begin
        IMAGE_addr <= 7976;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7999;
        test_state <= test_b1_S7993;
      end
      test_b1_S7993: begin
        IMAGE_addr <= 7977;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 583;
        test_state <= test_b1_S7994;
      end
      test_b1_S7994: begin
        IMAGE_addr <= 7978;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S7995;
      end
      test_b1_S7995: begin
        IMAGE_addr <= 7979;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5203;
        test_state <= test_b1_S7996;
      end
      test_b1_S7996: begin
        IMAGE_addr <= 7980;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S7997;
      end
      test_b1_S7997: begin
        IMAGE_addr <= 7981;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7995;
        test_state <= test_b1_S7998;
      end
      test_b1_S7998: begin
        IMAGE_addr <= 7982;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S7999;
      end
      test_b1_S7999: begin
        IMAGE_addr <= 7983;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7987;
        test_state <= test_b1_S8000;
      end
      test_b1_S8000: begin
        IMAGE_addr <= 7984;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 583;
        test_state <= test_b1_S8001;
      end
      test_b1_S8001: begin
        IMAGE_addr <= 7985;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S8002;
      end
      test_b1_S8002: begin
        IMAGE_addr <= 7986;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S8003;
      end
      test_b1_S8003: begin
        IMAGE_addr <= 7987;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S8004;
      end
      test_b1_S8004: begin
        IMAGE_addr <= 7988;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7992;
        test_state <= test_b1_S8005;
      end
      test_b1_S8005: begin
        IMAGE_addr <= 7989;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 578;
        test_state <= test_b1_S8006;
      end
      test_b1_S8006: begin
        IMAGE_addr <= 7990;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S8007;
      end
      test_b1_S8007: begin
        IMAGE_addr <= 7991;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S8008;
      end
      test_b1_S8008: begin
        IMAGE_addr <= 7992;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3539;
        test_state <= test_b1_S8009;
      end
      test_b1_S8009: begin
        IMAGE_addr <= 7993;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 183;
        test_state <= test_b1_S8010;
      end
      test_b1_S8010: begin
        IMAGE_addr <= 7994;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S8011;
      end
      test_b1_S8011: begin
        IMAGE_addr <= 7995;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S8012;
      end
      test_b1_S8012: begin
        IMAGE_addr <= 7996;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 52;
        test_state <= test_b1_S8013;
      end
      test_b1_S8013: begin
        IMAGE_addr <= 7997;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 732;
        test_state <= test_b1_S8014;
      end
      test_b1_S8014: begin
        IMAGE_addr <= 7998;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S8015;
      end
      test_b1_S8015: begin
        IMAGE_addr <= 7999;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S8016;
      end
      test_b1_S8016: begin
        IMAGE_addr <= 8000;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 52;
        test_state <= test_b1_S8017;
      end
      test_b1_S8017: begin
        IMAGE_addr <= 8001;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 732;
        test_state <= test_b1_S8018;
      end
      test_b1_S8018: begin
        IMAGE_addr <= 8002;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S8019;
      end
      test_b1_S8019: begin
        IMAGE_addr <= 8003;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S8020;
      end
      test_b1_S8020: begin
        IMAGE_addr <= 8004;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7962;
        test_state <= test_b1_S8021;
      end
      test_b1_S8021: begin
        IMAGE_addr <= 8005;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S8022;
      end
      test_b1_S8022: begin
        IMAGE_addr <= 8006;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8013;
        test_state <= test_b1_S8023;
      end
      test_b1_S8023: begin
        IMAGE_addr <= 8007;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 110;
        test_state <= test_b1_S8024;
      end
      test_b1_S8024: begin
        IMAGE_addr <= 8008;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S8025;
      end
      test_b1_S8025: begin
        IMAGE_addr <= 8009;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S8026;
      end
      test_b1_S8026: begin
        IMAGE_addr <= 8010;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 100;
        test_state <= test_b1_S8027;
      end
      test_b1_S8027: begin
        IMAGE_addr <= 8011;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S8028;
      end
      test_b1_S8028: begin
        IMAGE_addr <= 8012;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S8029;
      end
      test_b1_S8029: begin
        IMAGE_addr <= 8013;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S8030;
      end
      test_b1_S8030: begin
        IMAGE_addr <= 8014;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S8031;
      end
      test_b1_S8031: begin
        IMAGE_addr <= 8015;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6551;
        test_state <= test_b1_S8032;
      end
      test_b1_S8032: begin
        IMAGE_addr <= 8016;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S8033;
      end
      test_b1_S8033: begin
        IMAGE_addr <= 8017;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1232;
        test_state <= test_b1_S8034;
      end
      test_b1_S8034: begin
        IMAGE_addr <= 8018;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2577;
        test_state <= test_b1_S8035;
      end
      test_b1_S8035: begin
        IMAGE_addr <= 8019;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S8036;
      end
      test_b1_S8036: begin
        IMAGE_addr <= 8020;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 52;
        test_state <= test_b1_S8037;
      end
      test_b1_S8037: begin
        IMAGE_addr <= 8021;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S8038;
      end
      test_b1_S8038: begin
        IMAGE_addr <= 8022;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8049;
        test_state <= test_b1_S8039;
      end
      test_b1_S8039: begin
        IMAGE_addr <= 8023;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8;
        test_state <= test_b1_S8040;
      end
      test_b1_S8040: begin
        IMAGE_addr <= 8024;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8034;
        test_state <= test_b1_S8041;
      end
      test_b1_S8041: begin
        IMAGE_addr <= 8025;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 108;
        test_state <= test_b1_S8042;
      end
      test_b1_S8042: begin
        IMAGE_addr <= 8026;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S8043;
      end
      test_b1_S8043: begin
        IMAGE_addr <= 8027;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 98;
        test_state <= test_b1_S8044;
      end
      test_b1_S8044: begin
        IMAGE_addr <= 8028;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S8045;
      end
      test_b1_S8045: begin
        IMAGE_addr <= 8029;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S8046;
      end
      test_b1_S8046: begin
        IMAGE_addr <= 8030;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S8047;
      end
      test_b1_S8047: begin
        IMAGE_addr <= 8031;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 121;
        test_state <= test_b1_S8048;
      end
      test_b1_S8048: begin
        IMAGE_addr <= 8032;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 47;
        test_state <= test_b1_S8049;
      end
      test_b1_S8049: begin
        IMAGE_addr <= 8033;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S8050;
      end
      test_b1_S8050: begin
        IMAGE_addr <= 8034;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S8051;
      end
      test_b1_S8051: begin
        IMAGE_addr <= 8035;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8025;
        test_state <= test_b1_S8052;
      end
      test_b1_S8052: begin
        IMAGE_addr <= 8036;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7666;
        test_state <= test_b1_S8053;
      end
      test_b1_S8053: begin
        IMAGE_addr <= 8037;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7523;
        test_state <= test_b1_S8054;
      end
      test_b1_S8054: begin
        IMAGE_addr <= 8038;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8;
        test_state <= test_b1_S8055;
      end
      test_b1_S8055: begin
        IMAGE_addr <= 8039;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8044;
        test_state <= test_b1_S8056;
      end
      test_b1_S8056: begin
        IMAGE_addr <= 8040;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 46;
        test_state <= test_b1_S8057;
      end
      test_b1_S8057: begin
        IMAGE_addr <= 8041;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S8058;
      end
      test_b1_S8058: begin
        IMAGE_addr <= 8042;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 120;
        test_state <= test_b1_S8059;
      end
      test_b1_S8059: begin
        IMAGE_addr <= 8043;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S8060;
      end
      test_b1_S8060: begin
        IMAGE_addr <= 8044;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S8061;
      end
      test_b1_S8061: begin
        IMAGE_addr <= 8045;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8040;
        test_state <= test_b1_S8062;
      end
      test_b1_S8062: begin
        IMAGE_addr <= 8046;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 7700;
        test_state <= test_b1_S8063;
      end
      test_b1_S8063: begin
        IMAGE_addr <= 8047;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 6591;
        test_state <= test_b1_S8064;
      end
      test_b1_S8064: begin
        IMAGE_addr <= 8048;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S8065;
      end
      test_b1_S8065: begin
        IMAGE_addr <= 8049;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 732;
        test_state <= test_b1_S8066;
      end
      test_b1_S8066: begin
        IMAGE_addr <= 8050;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S8067;
      end
      test_b1_S8067: begin
        IMAGE_addr <= 8051;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S8068;
      end
      test_b1_S8068: begin
        IMAGE_addr <= 8052;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8004;
        test_state <= test_b1_S8069;
      end
      test_b1_S8069: begin
        IMAGE_addr <= 8053;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5034;
        test_state <= test_b1_S8070;
      end
      test_b1_S8070: begin
        IMAGE_addr <= 8054;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8426;
        test_state <= test_b1_S8071;
      end
      test_b1_S8071: begin
        IMAGE_addr <= 8055;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 102;
        test_state <= test_b1_S8072;
      end
      test_b1_S8072: begin
        IMAGE_addr <= 8056;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S8073;
      end
      test_b1_S8073: begin
        IMAGE_addr <= 8057;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 108;
        test_state <= test_b1_S8074;
      end
      test_b1_S8074: begin
        IMAGE_addr <= 8058;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S8075;
      end
      test_b1_S8075: begin
        IMAGE_addr <= 8059;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S8076;
      end
      test_b1_S8076: begin
        IMAGE_addr <= 8060;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 39;
        test_state <= test_b1_S8077;
      end
      test_b1_S8077: begin
        IMAGE_addr <= 8061;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S8078;
      end
      test_b1_S8078: begin
        IMAGE_addr <= 8062;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S8079;
      end
      test_b1_S8079: begin
        IMAGE_addr <= 8063;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S8080;
      end
      test_b1_S8080: begin
        IMAGE_addr <= 8064;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 306;
        test_state <= test_b1_S8081;
      end
      test_b1_S8081: begin
        IMAGE_addr <= 8065;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4956;
        test_state <= test_b1_S8082;
      end
      test_b1_S8082: begin
        IMAGE_addr <= 8066;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 37;
        test_state <= test_b1_S8083;
      end
      test_b1_S8083: begin
        IMAGE_addr <= 8067;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 37;
        test_state <= test_b1_S8084;
      end
      test_b1_S8084: begin
        IMAGE_addr <= 8068;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S8085;
      end
      test_b1_S8085: begin
        IMAGE_addr <= 8069;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8063;
        test_state <= test_b1_S8086;
      end
      test_b1_S8086: begin
        IMAGE_addr <= 8070;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 310;
        test_state <= test_b1_S8087;
      end
      test_b1_S8087: begin
        IMAGE_addr <= 8071;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8076;
        test_state <= test_b1_S8088;
      end
      test_b1_S8088: begin
        IMAGE_addr <= 8072;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 102;
        test_state <= test_b1_S8089;
      end
      test_b1_S8089: begin
        IMAGE_addr <= 8073;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S8090;
      end
      test_b1_S8090: begin
        IMAGE_addr <= 8074;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 100;
        test_state <= test_b1_S8091;
      end
      test_b1_S8091: begin
        IMAGE_addr <= 8075;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S8092;
      end
      test_b1_S8092: begin
        IMAGE_addr <= 8076;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S8093;
      end
      test_b1_S8093: begin
        IMAGE_addr <= 8077;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8069;
        test_state <= test_b1_S8094;
      end
      test_b1_S8094: begin
        IMAGE_addr <= 8078;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 310;
        test_state <= test_b1_S8095;
      end
      test_b1_S8095: begin
        IMAGE_addr <= 8079;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8086;
        test_state <= test_b1_S8096;
      end
      test_b1_S8096: begin
        IMAGE_addr <= 8080;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 102;
        test_state <= test_b1_S8097;
      end
      test_b1_S8097: begin
        IMAGE_addr <= 8081;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S8098;
      end
      test_b1_S8098: begin
        IMAGE_addr <= 8082;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S8099;
      end
      test_b1_S8099: begin
        IMAGE_addr <= 8083;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 122;
        test_state <= test_b1_S8100;
      end
      test_b1_S8100: begin
        IMAGE_addr <= 8084;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S8101;
      end
      test_b1_S8101: begin
        IMAGE_addr <= 8085;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S8102;
      end
      test_b1_S8102: begin
        IMAGE_addr <= 8086;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S8103;
      end
      test_b1_S8103: begin
        IMAGE_addr <= 8087;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8077;
        test_state <= test_b1_S8104;
      end
      test_b1_S8104: begin
        IMAGE_addr <= 8088;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 310;
        test_state <= test_b1_S8105;
      end
      test_b1_S8105: begin
        IMAGE_addr <= 8089;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8097;
        test_state <= test_b1_S8106;
      end
      test_b1_S8106: begin
        IMAGE_addr <= 8090;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S8107;
      end
      test_b1_S8107: begin
        IMAGE_addr <= 8091;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 99;
        test_state <= test_b1_S8108;
      end
      test_b1_S8108: begin
        IMAGE_addr <= 8092;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S8109;
      end
      test_b1_S8109: begin
        IMAGE_addr <= 8093;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S8110;
      end
      test_b1_S8110: begin
        IMAGE_addr <= 8094;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 118;
        test_state <= test_b1_S8111;
      end
      test_b1_S8111: begin
        IMAGE_addr <= 8095;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S8112;
      end
      test_b1_S8112: begin
        IMAGE_addr <= 8096;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S8113;
      end
      test_b1_S8113: begin
        IMAGE_addr <= 8097;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S8114;
      end
      test_b1_S8114: begin
        IMAGE_addr <= 8098;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8087;
        test_state <= test_b1_S8115;
      end
      test_b1_S8115: begin
        IMAGE_addr <= 8099;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S8116;
      end
      test_b1_S8116: begin
        IMAGE_addr <= 8100;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8104;
        test_state <= test_b1_S8117;
      end
      test_b1_S8117: begin
        IMAGE_addr <= 8101;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S8118;
      end
      test_b1_S8118: begin
        IMAGE_addr <= 8102;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 111;
        test_state <= test_b1_S8119;
      end
      test_b1_S8119: begin
        IMAGE_addr <= 8103;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S8120;
      end
      test_b1_S8120: begin
        IMAGE_addr <= 8104;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S8121;
      end
      test_b1_S8121: begin
        IMAGE_addr <= 8105;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S8122;
      end
      test_b1_S8122: begin
        IMAGE_addr <= 8106;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 29;
        test_state <= test_b1_S8123;
      end
      test_b1_S8123: begin
        IMAGE_addr <= 8107;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 122;
        test_state <= test_b1_S8124;
      end
      test_b1_S8124: begin
        IMAGE_addr <= 8108;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S8125;
      end
      test_b1_S8125: begin
        IMAGE_addr <= 8109;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S8126;
      end
      test_b1_S8126: begin
        IMAGE_addr <= 8110;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 28;
        test_state <= test_b1_S8127;
      end
      test_b1_S8127: begin
        IMAGE_addr <= 8111;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S8128;
      end
      test_b1_S8128: begin
        IMAGE_addr <= 8112;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S8129;
      end
      test_b1_S8129: begin
        IMAGE_addr <= 8113;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8098;
        test_state <= test_b1_S8130;
      end
      test_b1_S8130: begin
        IMAGE_addr <= 8114;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S8131;
      end
      test_b1_S8131: begin
        IMAGE_addr <= 8115;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8121;
        test_state <= test_b1_S8132;
      end
      test_b1_S8132: begin
        IMAGE_addr <= 8116;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 100;
        test_state <= test_b1_S8133;
      end
      test_b1_S8133: begin
        IMAGE_addr <= 8117;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 111;
        test_state <= test_b1_S8134;
      end
      test_b1_S8134: begin
        IMAGE_addr <= 8118;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 110;
        test_state <= test_b1_S8135;
      end
      test_b1_S8135: begin
        IMAGE_addr <= 8119;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S8136;
      end
      test_b1_S8136: begin
        IMAGE_addr <= 8120;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S8137;
      end
      test_b1_S8137: begin
        IMAGE_addr <= 8121;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S8138;
      end
      test_b1_S8138: begin
        IMAGE_addr <= 8122;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S8139;
      end
      test_b1_S8139: begin
        IMAGE_addr <= 8123;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S8140;
      end
      test_b1_S8140: begin
        IMAGE_addr <= 8124;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8097;
        test_state <= test_b1_S8141;
      end
      test_b1_S8141: begin
        IMAGE_addr <= 8125;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 155;
        test_state <= test_b1_S8142;
      end
      test_b1_S8142: begin
        IMAGE_addr <= 8126;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S8143;
      end
      test_b1_S8143: begin
        IMAGE_addr <= 8127;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S8144;
      end
      test_b1_S8144: begin
        IMAGE_addr <= 8128;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8063;
        test_state <= test_b1_S8145;
      end
      test_b1_S8145: begin
        IMAGE_addr <= 8129;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 310;
        test_state <= test_b1_S8146;
      end
      test_b1_S8146: begin
        IMAGE_addr <= 8130;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S8147;
      end
      test_b1_S8147: begin
        IMAGE_addr <= 8131;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 58;
        test_state <= test_b1_S8148;
      end
      test_b1_S8148: begin
        IMAGE_addr <= 8132;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 82;
        test_state <= test_b1_S8149;
      end
      test_b1_S8149: begin
        IMAGE_addr <= 8133;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S8150;
      end
      test_b1_S8150: begin
        IMAGE_addr <= 8134;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8128;
        test_state <= test_b1_S8151;
      end
      test_b1_S8151: begin
        IMAGE_addr <= 8135;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 310;
        test_state <= test_b1_S8152;
      end
      test_b1_S8152: begin
        IMAGE_addr <= 8136;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S8153;
      end
      test_b1_S8153: begin
        IMAGE_addr <= 8137;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 58;
        test_state <= test_b1_S8154;
      end
      test_b1_S8154: begin
        IMAGE_addr <= 8138;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 87;
        test_state <= test_b1_S8155;
      end
      test_b1_S8155: begin
        IMAGE_addr <= 8139;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S8156;
      end
      test_b1_S8156: begin
        IMAGE_addr <= 8140;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8134;
        test_state <= test_b1_S8157;
      end
      test_b1_S8157: begin
        IMAGE_addr <= 8141;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 310;
        test_state <= test_b1_S8158;
      end
      test_b1_S8158: begin
        IMAGE_addr <= 8142;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S8159;
      end
      test_b1_S8159: begin
        IMAGE_addr <= 8143;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 58;
        test_state <= test_b1_S8160;
      end
      test_b1_S8160: begin
        IMAGE_addr <= 8144;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 65;
        test_state <= test_b1_S8161;
      end
      test_b1_S8161: begin
        IMAGE_addr <= 8145;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S8162;
      end
      test_b1_S8162: begin
        IMAGE_addr <= 8146;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8140;
        test_state <= test_b1_S8163;
      end
      test_b1_S8163: begin
        IMAGE_addr <= 8147;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 310;
        test_state <= test_b1_S8164;
      end
      test_b1_S8164: begin
        IMAGE_addr <= 8148;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S8165;
      end
      test_b1_S8165: begin
        IMAGE_addr <= 8149;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 58;
        test_state <= test_b1_S8166;
      end
      test_b1_S8166: begin
        IMAGE_addr <= 8150;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 77;
        test_state <= test_b1_S8167;
      end
      test_b1_S8167: begin
        IMAGE_addr <= 8151;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S8168;
      end
      test_b1_S8168: begin
        IMAGE_addr <= 8152;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8146;
        test_state <= test_b1_S8169;
      end
      test_b1_S8169: begin
        IMAGE_addr <= 8153;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S8170;
      end
      test_b1_S8170: begin
        IMAGE_addr <= 8154;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8160;
        test_state <= test_b1_S8171;
      end
      test_b1_S8171: begin
        IMAGE_addr <= 8155;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 111;
        test_state <= test_b1_S8172;
      end
      test_b1_S8172: begin
        IMAGE_addr <= 8156;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 112;
        test_state <= test_b1_S8173;
      end
      test_b1_S8173: begin
        IMAGE_addr <= 8157;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S8174;
      end
      test_b1_S8174: begin
        IMAGE_addr <= 8158;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 110;
        test_state <= test_b1_S8175;
      end
      test_b1_S8175: begin
        IMAGE_addr <= 8159;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S8176;
      end
      test_b1_S8176: begin
        IMAGE_addr <= 8160;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S8177;
      end
      test_b1_S8177: begin
        IMAGE_addr <= 8161;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S8178;
      end
      test_b1_S8178: begin
        IMAGE_addr <= 8162;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S8179;
      end
      test_b1_S8179: begin
        IMAGE_addr <= 8163;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4294967295;
        test_state <= test_b1_S8180;
      end
      test_b1_S8180: begin
        IMAGE_addr <= 8164;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8104;
        test_state <= test_b1_S8181;
      end
      test_b1_S8181: begin
        IMAGE_addr <= 8165;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S8182;
      end
      test_b1_S8182: begin
        IMAGE_addr <= 8166;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S8183;
      end
      test_b1_S8183: begin
        IMAGE_addr <= 8167;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8152;
        test_state <= test_b1_S8184;
      end
      test_b1_S8184: begin
        IMAGE_addr <= 8168;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S8185;
      end
      test_b1_S8185: begin
        IMAGE_addr <= 8169;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8175;
        test_state <= test_b1_S8186;
      end
      test_b1_S8186: begin
        IMAGE_addr <= 8170;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S8187;
      end
      test_b1_S8187: begin
        IMAGE_addr <= 8171;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S8188;
      end
      test_b1_S8188: begin
        IMAGE_addr <= 8172;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S8189;
      end
      test_b1_S8189: begin
        IMAGE_addr <= 8173;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 100;
        test_state <= test_b1_S8190;
      end
      test_b1_S8190: begin
        IMAGE_addr <= 8174;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S8191;
      end
      test_b1_S8191: begin
        IMAGE_addr <= 8175;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S8192;
      end
      test_b1_S8192: begin
        IMAGE_addr <= 8176;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S8193;
      end
      test_b1_S8193: begin
        IMAGE_addr <= 8177;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S8194;
      end
      test_b1_S8194: begin
        IMAGE_addr <= 8178;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4294967294;
        test_state <= test_b1_S8195;
      end
      test_b1_S8195: begin
        IMAGE_addr <= 8179;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8104;
        test_state <= test_b1_S8196;
      end
      test_b1_S8196: begin
        IMAGE_addr <= 8180;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S8197;
      end
      test_b1_S8197: begin
        IMAGE_addr <= 8181;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S8198;
      end
      test_b1_S8198: begin
        IMAGE_addr <= 8182;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8167;
        test_state <= test_b1_S8199;
      end
      test_b1_S8199: begin
        IMAGE_addr <= 8183;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S8200;
      end
      test_b1_S8200: begin
        IMAGE_addr <= 8184;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8191;
        test_state <= test_b1_S8201;
      end
      test_b1_S8201: begin
        IMAGE_addr <= 8185;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 119;
        test_state <= test_b1_S8202;
      end
      test_b1_S8202: begin
        IMAGE_addr <= 8186;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S8203;
      end
      test_b1_S8203: begin
        IMAGE_addr <= 8187;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S8204;
      end
      test_b1_S8204: begin
        IMAGE_addr <= 8188;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S8205;
      end
      test_b1_S8205: begin
        IMAGE_addr <= 8189;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S8206;
      end
      test_b1_S8206: begin
        IMAGE_addr <= 8190;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S8207;
      end
      test_b1_S8207: begin
        IMAGE_addr <= 8191;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S8208;
      end
      test_b1_S8208: begin
        IMAGE_addr <= 8192;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S8209;
      end
      test_b1_S8209: begin
        IMAGE_addr <= 8193;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S8210;
      end
      test_b1_S8210: begin
        IMAGE_addr <= 8194;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4294967293;
        test_state <= test_b1_S8211;
      end
      test_b1_S8211: begin
        IMAGE_addr <= 8195;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8104;
        test_state <= test_b1_S8212;
      end
      test_b1_S8212: begin
        IMAGE_addr <= 8196;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S8213;
      end
      test_b1_S8213: begin
        IMAGE_addr <= 8197;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S8214;
      end
      test_b1_S8214: begin
        IMAGE_addr <= 8198;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8182;
        test_state <= test_b1_S8215;
      end
      test_b1_S8215: begin
        IMAGE_addr <= 8199;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S8216;
      end
      test_b1_S8216: begin
        IMAGE_addr <= 8200;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8207;
        test_state <= test_b1_S8217;
      end
      test_b1_S8217: begin
        IMAGE_addr <= 8201;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 99;
        test_state <= test_b1_S8218;
      end
      test_b1_S8218: begin
        IMAGE_addr <= 8202;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 108;
        test_state <= test_b1_S8219;
      end
      test_b1_S8219: begin
        IMAGE_addr <= 8203;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 111;
        test_state <= test_b1_S8220;
      end
      test_b1_S8220: begin
        IMAGE_addr <= 8204;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S8221;
      end
      test_b1_S8221: begin
        IMAGE_addr <= 8205;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S8222;
      end
      test_b1_S8222: begin
        IMAGE_addr <= 8206;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S8223;
      end
      test_b1_S8223: begin
        IMAGE_addr <= 8207;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S8224;
      end
      test_b1_S8224: begin
        IMAGE_addr <= 8208;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S8225;
      end
      test_b1_S8225: begin
        IMAGE_addr <= 8209;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S8226;
      end
      test_b1_S8226: begin
        IMAGE_addr <= 8210;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4294967292;
        test_state <= test_b1_S8227;
      end
      test_b1_S8227: begin
        IMAGE_addr <= 8211;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8104;
        test_state <= test_b1_S8228;
      end
      test_b1_S8228: begin
        IMAGE_addr <= 8212;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S8229;
      end
      test_b1_S8229: begin
        IMAGE_addr <= 8213;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S8230;
      end
      test_b1_S8230: begin
        IMAGE_addr <= 8214;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8198;
        test_state <= test_b1_S8231;
      end
      test_b1_S8231: begin
        IMAGE_addr <= 8215;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S8232;
      end
      test_b1_S8232: begin
        IMAGE_addr <= 8216;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8221;
        test_state <= test_b1_S8233;
      end
      test_b1_S8233: begin
        IMAGE_addr <= 8217;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 112;
        test_state <= test_b1_S8234;
      end
      test_b1_S8234: begin
        IMAGE_addr <= 8218;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 111;
        test_state <= test_b1_S8235;
      end
      test_b1_S8235: begin
        IMAGE_addr <= 8219;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S8236;
      end
      test_b1_S8236: begin
        IMAGE_addr <= 8220;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S8237;
      end
      test_b1_S8237: begin
        IMAGE_addr <= 8221;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S8238;
      end
      test_b1_S8238: begin
        IMAGE_addr <= 8222;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S8239;
      end
      test_b1_S8239: begin
        IMAGE_addr <= 8223;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S8240;
      end
      test_b1_S8240: begin
        IMAGE_addr <= 8224;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4294967291;
        test_state <= test_b1_S8241;
      end
      test_b1_S8241: begin
        IMAGE_addr <= 8225;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8104;
        test_state <= test_b1_S8242;
      end
      test_b1_S8242: begin
        IMAGE_addr <= 8226;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S8243;
      end
      test_b1_S8243: begin
        IMAGE_addr <= 8227;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S8244;
      end
      test_b1_S8244: begin
        IMAGE_addr <= 8228;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8214;
        test_state <= test_b1_S8245;
      end
      test_b1_S8245: begin
        IMAGE_addr <= 8229;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S8246;
      end
      test_b1_S8246: begin
        IMAGE_addr <= 8230;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8236;
        test_state <= test_b1_S8247;
      end
      test_b1_S8247: begin
        IMAGE_addr <= 8231;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S8248;
      end
      test_b1_S8248: begin
        IMAGE_addr <= 8232;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S8249;
      end
      test_b1_S8249: begin
        IMAGE_addr <= 8233;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S8250;
      end
      test_b1_S8250: begin
        IMAGE_addr <= 8234;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 107;
        test_state <= test_b1_S8251;
      end
      test_b1_S8251: begin
        IMAGE_addr <= 8235;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S8252;
      end
      test_b1_S8252: begin
        IMAGE_addr <= 8236;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S8253;
      end
      test_b1_S8253: begin
        IMAGE_addr <= 8237;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S8254;
      end
      test_b1_S8254: begin
        IMAGE_addr <= 8238;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S8255;
      end
      test_b1_S8255: begin
        IMAGE_addr <= 8239;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4294967290;
        test_state <= test_b1_S8256;
      end
      test_b1_S8256: begin
        IMAGE_addr <= 8240;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8104;
        test_state <= test_b1_S8257;
      end
      test_b1_S8257: begin
        IMAGE_addr <= 8241;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S8258;
      end
      test_b1_S8258: begin
        IMAGE_addr <= 8242;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S8259;
      end
      test_b1_S8259: begin
        IMAGE_addr <= 8243;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8228;
        test_state <= test_b1_S8260;
      end
      test_b1_S8260: begin
        IMAGE_addr <= 8244;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S8261;
      end
      test_b1_S8261: begin
        IMAGE_addr <= 8245;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8251;
        test_state <= test_b1_S8262;
      end
      test_b1_S8262: begin
        IMAGE_addr <= 8246;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S8263;
      end
      test_b1_S8263: begin
        IMAGE_addr <= 8247;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S8264;
      end
      test_b1_S8264: begin
        IMAGE_addr <= 8248;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 122;
        test_state <= test_b1_S8265;
      end
      test_b1_S8265: begin
        IMAGE_addr <= 8249;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S8266;
      end
      test_b1_S8266: begin
        IMAGE_addr <= 8250;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S8267;
      end
      test_b1_S8267: begin
        IMAGE_addr <= 8251;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S8268;
      end
      test_b1_S8268: begin
        IMAGE_addr <= 8252;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S8269;
      end
      test_b1_S8269: begin
        IMAGE_addr <= 8253;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S8270;
      end
      test_b1_S8270: begin
        IMAGE_addr <= 8254;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4294967289;
        test_state <= test_b1_S8271;
      end
      test_b1_S8271: begin
        IMAGE_addr <= 8255;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8104;
        test_state <= test_b1_S8272;
      end
      test_b1_S8272: begin
        IMAGE_addr <= 8256;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S8273;
      end
      test_b1_S8273: begin
        IMAGE_addr <= 8257;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S8274;
      end
      test_b1_S8274: begin
        IMAGE_addr <= 8258;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8243;
        test_state <= test_b1_S8275;
      end
      test_b1_S8275: begin
        IMAGE_addr <= 8259;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S8276;
      end
      test_b1_S8276: begin
        IMAGE_addr <= 8260;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8268;
        test_state <= test_b1_S8277;
      end
      test_b1_S8277: begin
        IMAGE_addr <= 8261;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 100;
        test_state <= test_b1_S8278;
      end
      test_b1_S8278: begin
        IMAGE_addr <= 8262;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S8279;
      end
      test_b1_S8279: begin
        IMAGE_addr <= 8263;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 108;
        test_state <= test_b1_S8280;
      end
      test_b1_S8280: begin
        IMAGE_addr <= 8264;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S8281;
      end
      test_b1_S8281: begin
        IMAGE_addr <= 8265;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S8282;
      end
      test_b1_S8282: begin
        IMAGE_addr <= 8266;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S8283;
      end
      test_b1_S8283: begin
        IMAGE_addr <= 8267;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S8284;
      end
      test_b1_S8284: begin
        IMAGE_addr <= 8268;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S8285;
      end
      test_b1_S8285: begin
        IMAGE_addr <= 8269;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S8286;
      end
      test_b1_S8286: begin
        IMAGE_addr <= 8270;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S8287;
      end
      test_b1_S8287: begin
        IMAGE_addr <= 8271;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4294967288;
        test_state <= test_b1_S8288;
      end
      test_b1_S8288: begin
        IMAGE_addr <= 8272;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8104;
        test_state <= test_b1_S8289;
      end
      test_b1_S8289: begin
        IMAGE_addr <= 8273;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S8290;
      end
      test_b1_S8290: begin
        IMAGE_addr <= 8274;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S8291;
      end
      test_b1_S8291: begin
        IMAGE_addr <= 8275;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8258;
        test_state <= test_b1_S8292;
      end
      test_b1_S8292: begin
        IMAGE_addr <= 8276;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S8293;
      end
      test_b1_S8293: begin
        IMAGE_addr <= 8277;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8284;
        test_state <= test_b1_S8294;
      end
      test_b1_S8294: begin
        IMAGE_addr <= 8278;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S8295;
      end
      test_b1_S8295: begin
        IMAGE_addr <= 8279;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 108;
        test_state <= test_b1_S8296;
      end
      test_b1_S8296: begin
        IMAGE_addr <= 8280;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 117;
        test_state <= test_b1_S8297;
      end
      test_b1_S8297: begin
        IMAGE_addr <= 8281;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S8298;
      end
      test_b1_S8298: begin
        IMAGE_addr <= 8282;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 112;
        test_state <= test_b1_S8299;
      end
      test_b1_S8299: begin
        IMAGE_addr <= 8283;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S8300;
      end
      test_b1_S8300: begin
        IMAGE_addr <= 8284;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S8301;
      end
      test_b1_S8301: begin
        IMAGE_addr <= 8285;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S8302;
      end
      test_b1_S8302: begin
        IMAGE_addr <= 8286;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S8303;
      end
      test_b1_S8303: begin
        IMAGE_addr <= 8287;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S8304;
      end
      test_b1_S8304: begin
        IMAGE_addr <= 8288;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8160;
        test_state <= test_b1_S8305;
      end
      test_b1_S8305: begin
        IMAGE_addr <= 8289;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S8306;
      end
      test_b1_S8306: begin
        IMAGE_addr <= 8290;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8076;
        test_state <= test_b1_S8307;
      end
      test_b1_S8307: begin
        IMAGE_addr <= 8291;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S8308;
      end
      test_b1_S8308: begin
        IMAGE_addr <= 8292;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S8309;
      end
      test_b1_S8309: begin
        IMAGE_addr <= 8293;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8076;
        test_state <= test_b1_S8310;
      end
      test_b1_S8310: begin
        IMAGE_addr <= 8294;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S8311;
      end
      test_b1_S8311: begin
        IMAGE_addr <= 8295;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8251;
        test_state <= test_b1_S8312;
      end
      test_b1_S8312: begin
        IMAGE_addr <= 8296;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S8313;
      end
      test_b1_S8313: begin
        IMAGE_addr <= 8297;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8086;
        test_state <= test_b1_S8314;
      end
      test_b1_S8314: begin
        IMAGE_addr <= 8298;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S8315;
      end
      test_b1_S8315: begin
        IMAGE_addr <= 8299;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S8316;
      end
      test_b1_S8316: begin
        IMAGE_addr <= 8300;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8086;
        test_state <= test_b1_S8317;
      end
      test_b1_S8317: begin
        IMAGE_addr <= 8301;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S8318;
      end
      test_b1_S8318: begin
        IMAGE_addr <= 8302;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S8319;
      end
      test_b1_S8319: begin
        IMAGE_addr <= 8303;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8311;
        test_state <= test_b1_S8320;
      end
      test_b1_S8320: begin
        IMAGE_addr <= 8304;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S8321;
      end
      test_b1_S8321: begin
        IMAGE_addr <= 8305;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8076;
        test_state <= test_b1_S8322;
      end
      test_b1_S8322: begin
        IMAGE_addr <= 8306;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S8323;
      end
      test_b1_S8323: begin
        IMAGE_addr <= 8307;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8175;
        test_state <= test_b1_S8324;
      end
      test_b1_S8324: begin
        IMAGE_addr <= 8308;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S8325;
      end
      test_b1_S8325: begin
        IMAGE_addr <= 8309;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 197;
        test_state <= test_b1_S8326;
      end
      test_b1_S8326: begin
        IMAGE_addr <= 8310;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S8327;
      end
      test_b1_S8327: begin
        IMAGE_addr <= 8311;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3841;
        test_state <= test_b1_S8328;
      end
      test_b1_S8328: begin
        IMAGE_addr <= 8312;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S8329;
      end
      test_b1_S8329: begin
        IMAGE_addr <= 8313;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S8330;
      end
      test_b1_S8330: begin
        IMAGE_addr <= 8314;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S8331;
      end
      test_b1_S8331: begin
        IMAGE_addr <= 8315;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S8332;
      end
      test_b1_S8332: begin
        IMAGE_addr <= 8316;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S8333;
      end
      test_b1_S8333: begin
        IMAGE_addr <= 8317;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8076;
        test_state <= test_b1_S8334;
      end
      test_b1_S8334: begin
        IMAGE_addr <= 8318;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S8335;
      end
      test_b1_S8335: begin
        IMAGE_addr <= 8319;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8207;
        test_state <= test_b1_S8336;
      end
      test_b1_S8336: begin
        IMAGE_addr <= 8320;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S8337;
      end
      test_b1_S8337: begin
        IMAGE_addr <= 8321;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S8338;
      end
      test_b1_S8338: begin
        IMAGE_addr <= 8322;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8086;
        test_state <= test_b1_S8339;
      end
      test_b1_S8339: begin
        IMAGE_addr <= 8323;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S8340;
      end
      test_b1_S8340: begin
        IMAGE_addr <= 8324;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S8341;
      end
      test_b1_S8341: begin
        IMAGE_addr <= 8325;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S8342;
      end
      test_b1_S8342: begin
        IMAGE_addr <= 8326;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8275;
        test_state <= test_b1_S8343;
      end
      test_b1_S8343: begin
        IMAGE_addr <= 8327;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S8344;
      end
      test_b1_S8344: begin
        IMAGE_addr <= 8328;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8334;
        test_state <= test_b1_S8345;
      end
      test_b1_S8345: begin
        IMAGE_addr <= 8329;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S8346;
      end
      test_b1_S8346: begin
        IMAGE_addr <= 8330;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 112;
        test_state <= test_b1_S8347;
      end
      test_b1_S8347: begin
        IMAGE_addr <= 8331;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S8348;
      end
      test_b1_S8348: begin
        IMAGE_addr <= 8332;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 119;
        test_state <= test_b1_S8349;
      end
      test_b1_S8349: begin
        IMAGE_addr <= 8333;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S8350;
      end
      test_b1_S8350: begin
        IMAGE_addr <= 8334;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S8351;
      end
      test_b1_S8351: begin
        IMAGE_addr <= 8335;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S8352;
      end
      test_b1_S8352: begin
        IMAGE_addr <= 8336;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S8353;
      end
      test_b1_S8353: begin
        IMAGE_addr <= 8337;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S8354;
      end
      test_b1_S8354: begin
        IMAGE_addr <= 8338;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8160;
        test_state <= test_b1_S8355;
      end
      test_b1_S8355: begin
        IMAGE_addr <= 8339;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S8356;
      end
      test_b1_S8356: begin
        IMAGE_addr <= 8340;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8076;
        test_state <= test_b1_S8357;
      end
      test_b1_S8357: begin
        IMAGE_addr <= 8341;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S8358;
      end
      test_b1_S8358: begin
        IMAGE_addr <= 8342;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S8359;
      end
      test_b1_S8359: begin
        IMAGE_addr <= 8343;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S8360;
      end
      test_b1_S8360: begin
        IMAGE_addr <= 8344;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S8361;
      end
      test_b1_S8361: begin
        IMAGE_addr <= 8345;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8086;
        test_state <= test_b1_S8362;
      end
      test_b1_S8362: begin
        IMAGE_addr <= 8346;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S8363;
      end
      test_b1_S8363: begin
        IMAGE_addr <= 8347;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S8364;
      end
      test_b1_S8364: begin
        IMAGE_addr <= 8348;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8359;
        test_state <= test_b1_S8365;
      end
      test_b1_S8365: begin
        IMAGE_addr <= 8349;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 189;
        test_state <= test_b1_S8366;
      end
      test_b1_S8366: begin
        IMAGE_addr <= 8350;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S8367;
      end
      test_b1_S8367: begin
        IMAGE_addr <= 8351;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8076;
        test_state <= test_b1_S8368;
      end
      test_b1_S8368: begin
        IMAGE_addr <= 8352;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S8369;
      end
      test_b1_S8369: begin
        IMAGE_addr <= 8353;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8191;
        test_state <= test_b1_S8370;
      end
      test_b1_S8370: begin
        IMAGE_addr <= 8354;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S8371;
      end
      test_b1_S8371: begin
        IMAGE_addr <= 8355;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S8372;
      end
      test_b1_S8372: begin
        IMAGE_addr <= 8356;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8086;
        test_state <= test_b1_S8373;
      end
      test_b1_S8373: begin
        IMAGE_addr <= 8357;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2651;
        test_state <= test_b1_S8374;
      end
      test_b1_S8374: begin
        IMAGE_addr <= 8358;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S8375;
      end
      test_b1_S8375: begin
        IMAGE_addr <= 8359;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3841;
        test_state <= test_b1_S8376;
      end
      test_b1_S8376: begin
        IMAGE_addr <= 8360;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S8377;
      end
      test_b1_S8377: begin
        IMAGE_addr <= 8361;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S8378;
      end
      test_b1_S8378: begin
        IMAGE_addr <= 8362;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8076;
        test_state <= test_b1_S8379;
      end
      test_b1_S8379: begin
        IMAGE_addr <= 8363;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S8380;
      end
      test_b1_S8380: begin
        IMAGE_addr <= 8364;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8207;
        test_state <= test_b1_S8381;
      end
      test_b1_S8381: begin
        IMAGE_addr <= 8365;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S8382;
      end
      test_b1_S8382: begin
        IMAGE_addr <= 8366;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S8383;
      end
      test_b1_S8383: begin
        IMAGE_addr <= 8367;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8086;
        test_state <= test_b1_S8384;
      end
      test_b1_S8384: begin
        IMAGE_addr <= 8368;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S8385;
      end
      test_b1_S8385: begin
        IMAGE_addr <= 8369;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S8386;
      end
      test_b1_S8386: begin
        IMAGE_addr <= 8370;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S8387;
      end
      test_b1_S8387: begin
        IMAGE_addr <= 8371;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8326;
        test_state <= test_b1_S8388;
      end
      test_b1_S8388: begin
        IMAGE_addr <= 8372;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S8389;
      end
      test_b1_S8389: begin
        IMAGE_addr <= 8373;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8383;
        test_state <= test_b1_S8390;
      end
      test_b1_S8390: begin
        IMAGE_addr <= 8374;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S8391;
      end
      test_b1_S8391: begin
        IMAGE_addr <= 8375;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S8392;
      end
      test_b1_S8392: begin
        IMAGE_addr <= 8376;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 97;
        test_state <= test_b1_S8393;
      end
      test_b1_S8393: begin
        IMAGE_addr <= 8377;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 100;
        test_state <= test_b1_S8394;
      end
      test_b1_S8394: begin
        IMAGE_addr <= 8378;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 76;
        test_state <= test_b1_S8395;
      end
      test_b1_S8395: begin
        IMAGE_addr <= 8379;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S8396;
      end
      test_b1_S8396: begin
        IMAGE_addr <= 8380;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 110;
        test_state <= test_b1_S8397;
      end
      test_b1_S8397: begin
        IMAGE_addr <= 8381;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S8398;
      end
      test_b1_S8398: begin
        IMAGE_addr <= 8382;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S8399;
      end
      test_b1_S8399: begin
        IMAGE_addr <= 8383;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S8400;
      end
      test_b1_S8400: begin
        IMAGE_addr <= 8384;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S8401;
      end
      test_b1_S8401: begin
        IMAGE_addr <= 8385;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S8402;
      end
      test_b1_S8402: begin
        IMAGE_addr <= 8386;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8097;
        test_state <= test_b1_S8403;
      end
      test_b1_S8403: begin
        IMAGE_addr <= 8387;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 147;
        test_state <= test_b1_S8404;
      end
      test_b1_S8404: begin
        IMAGE_addr <= 8388;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 400;
        test_state <= test_b1_S8405;
      end
      test_b1_S8405: begin
        IMAGE_addr <= 8389;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S8406;
      end
      test_b1_S8406: begin
        IMAGE_addr <= 8390;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8421;
        test_state <= test_b1_S8407;
      end
      test_b1_S8407: begin
        IMAGE_addr <= 8391;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 132;
        test_state <= test_b1_S8408;
      end
      test_b1_S8408: begin
        IMAGE_addr <= 8392;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8175;
        test_state <= test_b1_S8409;
      end
      test_b1_S8409: begin
        IMAGE_addr <= 8393;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S8410;
      end
      test_b1_S8410: begin
        IMAGE_addr <= 8394;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S8411;
      end
      test_b1_S8411: begin
        IMAGE_addr <= 8395;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 10;
        test_state <= test_b1_S8412;
      end
      test_b1_S8412: begin
        IMAGE_addr <= 8396;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S8413;
      end
      test_b1_S8413: begin
        IMAGE_addr <= 8397;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 13;
        test_state <= test_b1_S8414;
      end
      test_b1_S8414: begin
        IMAGE_addr <= 8398;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4214;
        test_state <= test_b1_S8415;
      end
      test_b1_S8415: begin
        IMAGE_addr <= 8399;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S8416;
      end
      test_b1_S8416: begin
        IMAGE_addr <= 8400;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8411;
        test_state <= test_b1_S8417;
      end
      test_b1_S8417: begin
        IMAGE_addr <= 8401;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S8418;
      end
      test_b1_S8418: begin
        IMAGE_addr <= 8402;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S8419;
      end
      test_b1_S8419: begin
        IMAGE_addr <= 8403;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S8420;
      end
      test_b1_S8420: begin
        IMAGE_addr <= 8404;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S8421;
      end
      test_b1_S8421: begin
        IMAGE_addr <= 8405;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S8422;
      end
      test_b1_S8422: begin
        IMAGE_addr <= 8406;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S8423;
      end
      test_b1_S8423: begin
        IMAGE_addr <= 8407;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S8424;
      end
      test_b1_S8424: begin
        IMAGE_addr <= 8408;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8097;
        test_state <= test_b1_S8425;
      end
      test_b1_S8425: begin
        IMAGE_addr <= 8409;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 155;
        test_state <= test_b1_S8426;
      end
      test_b1_S8426: begin
        IMAGE_addr <= 8410;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S8427;
      end
      test_b1_S8427: begin
        IMAGE_addr <= 8411;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S8428;
      end
      test_b1_S8428: begin
        IMAGE_addr <= 8412;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8416;
        test_state <= test_b1_S8429;
      end
      test_b1_S8429: begin
        IMAGE_addr <= 8413;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4;
        test_state <= test_b1_S8430;
      end
      test_b1_S8430: begin
        IMAGE_addr <= 8414;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 197;
        test_state <= test_b1_S8431;
      end
      test_b1_S8431: begin
        IMAGE_addr <= 8415;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S8432;
      end
      test_b1_S8432: begin
        IMAGE_addr <= 8416;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 732;
        test_state <= test_b1_S8433;
      end
      test_b1_S8433: begin
        IMAGE_addr <= 8417;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S8434;
      end
      test_b1_S8434: begin
        IMAGE_addr <= 8418;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8097;
        test_state <= test_b1_S8435;
      end
      test_b1_S8435: begin
        IMAGE_addr <= 8419;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S8436;
      end
      test_b1_S8436: begin
        IMAGE_addr <= 8420;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S8437;
      end
      test_b1_S8437: begin
        IMAGE_addr <= 8421;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3433;
        test_state <= test_b1_S8438;
      end
      test_b1_S8438: begin
        IMAGE_addr <= 8422;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 400;
        test_state <= test_b1_S8439;
      end
      test_b1_S8439: begin
        IMAGE_addr <= 8423;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5792;
        test_state <= test_b1_S8440;
      end
      test_b1_S8440: begin
        IMAGE_addr <= 8424;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S8441;
      end
      test_b1_S8441: begin
        IMAGE_addr <= 8425;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S8442;
      end
      test_b1_S8442: begin
        IMAGE_addr <= 8426;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8371;
        test_state <= test_b1_S8443;
      end
      test_b1_S8443: begin
        IMAGE_addr <= 8427;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 292;
        test_state <= test_b1_S8444;
      end
      test_b1_S8444: begin
        IMAGE_addr <= 8428;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8439;
        test_state <= test_b1_S8445;
      end
      test_b1_S8445: begin
        IMAGE_addr <= 8429;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 119;
        test_state <= test_b1_S8446;
      end
      test_b1_S8446: begin
        IMAGE_addr <= 8430;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 114;
        test_state <= test_b1_S8447;
      end
      test_b1_S8447: begin
        IMAGE_addr <= 8431;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S8448;
      end
      test_b1_S8448: begin
        IMAGE_addr <= 8432;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S8449;
      end
      test_b1_S8449: begin
        IMAGE_addr <= 8433;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S8450;
      end
      test_b1_S8450: begin
        IMAGE_addr <= 8434;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 76;
        test_state <= test_b1_S8451;
      end
      test_b1_S8451: begin
        IMAGE_addr <= 8435;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 105;
        test_state <= test_b1_S8452;
      end
      test_b1_S8452: begin
        IMAGE_addr <= 8436;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 110;
        test_state <= test_b1_S8453;
      end
      test_b1_S8453: begin
        IMAGE_addr <= 8437;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S8454;
      end
      test_b1_S8454: begin
        IMAGE_addr <= 8438;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S8455;
      end
      test_b1_S8455: begin
        IMAGE_addr <= 8439;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S8456;
      end
      test_b1_S8456: begin
        IMAGE_addr <= 8440;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S8457;
      end
      test_b1_S8457: begin
        IMAGE_addr <= 8441;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S8458;
      end
      test_b1_S8458: begin
        IMAGE_addr <= 8442;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8076;
        test_state <= test_b1_S8459;
      end
      test_b1_S8459: begin
        IMAGE_addr <= 8443;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 15;
        test_state <= test_b1_S8460;
      end
      test_b1_S8460: begin
        IMAGE_addr <= 8444;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S8461;
      end
      test_b1_S8461: begin
        IMAGE_addr <= 8445;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8097;
        test_state <= test_b1_S8462;
      end
      test_b1_S8462: begin
        IMAGE_addr <= 8446;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 147;
        test_state <= test_b1_S8463;
      end
      test_b1_S8463: begin
        IMAGE_addr <= 8447;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S8464;
      end
      test_b1_S8464: begin
        IMAGE_addr <= 8448;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8469;
        test_state <= test_b1_S8465;
      end
      test_b1_S8465: begin
        IMAGE_addr <= 8449;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 189;
        test_state <= test_b1_S8466;
      end
      test_b1_S8466: begin
        IMAGE_addr <= 8450;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S8467;
      end
      test_b1_S8467: begin
        IMAGE_addr <= 8451;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S8468;
      end
      test_b1_S8468: begin
        IMAGE_addr <= 8452;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S8469;
      end
      test_b1_S8469: begin
        IMAGE_addr <= 8453;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 790;
        test_state <= test_b1_S8470;
      end
      test_b1_S8470: begin
        IMAGE_addr <= 8454;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S8471;
      end
      test_b1_S8471: begin
        IMAGE_addr <= 8455;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8121;
        test_state <= test_b1_S8472;
      end
      test_b1_S8472: begin
        IMAGE_addr <= 8456;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 680;
        test_state <= test_b1_S8473;
      end
      test_b1_S8473: begin
        IMAGE_addr <= 8457;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8464;
        test_state <= test_b1_S8474;
      end
      test_b1_S8474: begin
        IMAGE_addr <= 8458;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S8475;
      end
      test_b1_S8475: begin
        IMAGE_addr <= 8459;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8076;
        test_state <= test_b1_S8476;
      end
      test_b1_S8476: begin
        IMAGE_addr <= 8460;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S8477;
      end
      test_b1_S8477: begin
        IMAGE_addr <= 8461;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8191;
        test_state <= test_b1_S8478;
      end
      test_b1_S8478: begin
        IMAGE_addr <= 8462;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S8479;
      end
      test_b1_S8479: begin
        IMAGE_addr <= 8463;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S8480;
      end
      test_b1_S8480: begin
        IMAGE_addr <= 8464;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 732;
        test_state <= test_b1_S8481;
      end
      test_b1_S8481: begin
        IMAGE_addr <= 8465;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S8482;
      end
      test_b1_S8482: begin
        IMAGE_addr <= 8466;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8097;
        test_state <= test_b1_S8483;
      end
      test_b1_S8483: begin
        IMAGE_addr <= 8467;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S8484;
      end
      test_b1_S8484: begin
        IMAGE_addr <= 8468;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S8485;
      end
      test_b1_S8485: begin
        IMAGE_addr <= 8469;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3433;
        test_state <= test_b1_S8486;
      end
      test_b1_S8486: begin
        IMAGE_addr <= 8470;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S8487;
      end
      test_b1_S8487: begin
        IMAGE_addr <= 8471;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 10;
        test_state <= test_b1_S8488;
      end
      test_b1_S8488: begin
        IMAGE_addr <= 8472;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S8489;
      end
      test_b1_S8489: begin
        IMAGE_addr <= 8473;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8076;
        test_state <= test_b1_S8490;
      end
      test_b1_S8490: begin
        IMAGE_addr <= 8474;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 14;
        test_state <= test_b1_S8491;
      end
      test_b1_S8491: begin
        IMAGE_addr <= 8475;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8191;
        test_state <= test_b1_S8492;
      end
      test_b1_S8492: begin
        IMAGE_addr <= 8476;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S8493;
      end
      test_b1_S8493: begin
        IMAGE_addr <= 8477;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S8494;
      end
      test_b1_S8494: begin
        IMAGE_addr <= 8478;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 9;
        test_state <= test_b1_S8495;
      end
      test_b1_S8495: begin
        IMAGE_addr <= 8479;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8052;
        test_state <= test_b1_S8496;
      end
      test_b1_S8496: begin
        IMAGE_addr <= 8480;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 5034;
        test_state <= test_b1_S8497;
      end
      test_b1_S8497: begin
        IMAGE_addr <= 8481;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8525;
        test_state <= test_b1_S8498;
      end
      test_b1_S8498: begin
        IMAGE_addr <= 8482;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 116;
        test_state <= test_b1_S8499;
      end
      test_b1_S8499: begin
        IMAGE_addr <= 8483;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 121;
        test_state <= test_b1_S8500;
      end
      test_b1_S8500: begin
        IMAGE_addr <= 8484;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 112;
        test_state <= test_b1_S8501;
      end
      test_b1_S8501: begin
        IMAGE_addr <= 8485;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 101;
        test_state <= test_b1_S8502;
      end
      test_b1_S8502: begin
        IMAGE_addr <= 8486;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 115;
        test_state <= test_b1_S8503;
      end
      test_b1_S8503: begin
        IMAGE_addr <= 8487;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 39;
        test_state <= test_b1_S8504;
      end
      test_b1_S8504: begin
        IMAGE_addr <= 8488;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S8505;
      end
      test_b1_S8505: begin
        IMAGE_addr <= 8489;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S8506;
      end
      test_b1_S8506: begin
        IMAGE_addr <= 8490;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S8507;
      end
      test_b1_S8507: begin
        IMAGE_addr <= 8491;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 306;
        test_state <= test_b1_S8508;
      end
      test_b1_S8508: begin
        IMAGE_addr <= 8492;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 4956;
        test_state <= test_b1_S8509;
      end
      test_b1_S8509: begin
        IMAGE_addr <= 8493;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 37;
        test_state <= test_b1_S8510;
      end
      test_b1_S8510: begin
        IMAGE_addr <= 8494;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 37;
        test_state <= test_b1_S8511;
      end
      test_b1_S8511: begin
        IMAGE_addr <= 8495;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S8512;
      end
      test_b1_S8512: begin
        IMAGE_addr <= 8496;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8490;
        test_state <= test_b1_S8513;
      end
      test_b1_S8513: begin
        IMAGE_addr <= 8497;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 310;
        test_state <= test_b1_S8514;
      end
      test_b1_S8514: begin
        IMAGE_addr <= 8498;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S8515;
      end
      test_b1_S8515: begin
        IMAGE_addr <= 8499;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 65;
        test_state <= test_b1_S8516;
      end
      test_b1_S8516: begin
        IMAGE_addr <= 8500;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 82;
        test_state <= test_b1_S8517;
      end
      test_b1_S8517: begin
        IMAGE_addr <= 8501;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 82;
        test_state <= test_b1_S8518;
      end
      test_b1_S8518: begin
        IMAGE_addr <= 8502;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 65;
        test_state <= test_b1_S8519;
      end
      test_b1_S8519: begin
        IMAGE_addr <= 8503;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 89;
        test_state <= test_b1_S8520;
      end
      test_b1_S8520: begin
        IMAGE_addr <= 8504;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S8521;
      end
      test_b1_S8521: begin
        IMAGE_addr <= 8505;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8496;
        test_state <= test_b1_S8522;
      end
      test_b1_S8522: begin
        IMAGE_addr <= 8506;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 310;
        test_state <= test_b1_S8523;
      end
      test_b1_S8523: begin
        IMAGE_addr <= 8507;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 1;
        test_state <= test_b1_S8524;
      end
      test_b1_S8524: begin
        IMAGE_addr <= 8508;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 66;
        test_state <= test_b1_S8525;
      end
      test_b1_S8525: begin
        IMAGE_addr <= 8509;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 85;
        test_state <= test_b1_S8526;
      end
      test_b1_S8526: begin
        IMAGE_addr <= 8510;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 70;
        test_state <= test_b1_S8527;
      end
      test_b1_S8527: begin
        IMAGE_addr <= 8511;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 70;
        test_state <= test_b1_S8528;
      end
      test_b1_S8528: begin
        IMAGE_addr <= 8512;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 69;
        test_state <= test_b1_S8529;
      end
      test_b1_S8529: begin
        IMAGE_addr <= 8513;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 82;
        test_state <= test_b1_S8530;
      end
      test_b1_S8530: begin
        IMAGE_addr <= 8514;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S8531;
      end
      test_b1_S8531: begin
        IMAGE_addr <= 8515;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8505;
        test_state <= test_b1_S8532;
      end
      test_b1_S8532: begin
        IMAGE_addr <= 8516;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 310;
        test_state <= test_b1_S8533;
      end
      test_b1_S8533: begin
        IMAGE_addr <= 8517;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 2;
        test_state <= test_b1_S8534;
      end
      test_b1_S8534: begin
        IMAGE_addr <= 8518;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 83;
        test_state <= test_b1_S8535;
      end
      test_b1_S8535: begin
        IMAGE_addr <= 8519;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 84;
        test_state <= test_b1_S8536;
      end
      test_b1_S8536: begin
        IMAGE_addr <= 8520;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 82;
        test_state <= test_b1_S8537;
      end
      test_b1_S8537: begin
        IMAGE_addr <= 8521;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 73;
        test_state <= test_b1_S8538;
      end
      test_b1_S8538: begin
        IMAGE_addr <= 8522;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 78;
        test_state <= test_b1_S8539;
      end
      test_b1_S8539: begin
        IMAGE_addr <= 8523;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 71;
        test_state <= test_b1_S8540;
      end
      test_b1_S8540: begin
        IMAGE_addr <= 8524;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S8541;
      end
      test_b1_S8541: begin
        IMAGE_addr <= 8525;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 8515;
        test_state <= test_b1_S8542;
      end
      test_b1_S8542: begin
        IMAGE_addr <= 8526;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 310;
        test_state <= test_b1_S8543;
      end
      test_b1_S8543: begin
        IMAGE_addr <= 8527;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 3;
        test_state <= test_b1_S8544;
      end
      test_b1_S8544: begin
        IMAGE_addr <= 8528;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 76;
        test_state <= test_b1_S8545;
      end
      test_b1_S8545: begin
        IMAGE_addr <= 8529;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 73;
        test_state <= test_b1_S8546;
      end
      test_b1_S8546: begin
        IMAGE_addr <= 8530;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 83;
        test_state <= test_b1_S8547;
      end
      test_b1_S8547: begin
        IMAGE_addr <= 8531;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 84;
        test_state <= test_b1_S8548;
      end
      test_b1_S8548: begin
        IMAGE_addr <= 8532;
        IMAGE_we <= 1;
        IMAGE_req <= 1;
        IMAGE_d <= 0;
        test_state <= test_b1_S8549;
      end
      test_b1_S8549: begin
        retro_main_0_ready <= 1;
        IMAGE_req <= 0;
        test_state <= test_b1_S8550;
      end
      test_b1_S8550: begin
        retro_main_0_ready <= 0;
        test_state <= test_b1_S8551;
      end
      test_b1_S8551: begin
        if (retro_main_0_valid == 1) begin
          retro_main_0_accept <= 1;
          test_state <= test_b1_S8553;
        end
      end
      test_b1_S8553: begin
        retro_main_0_accept <= 0;
        test_state <= test_b1_FINISH;
      end
      test_b1_FINISH: begin
        $display("%5t:finish", $time);
        $finish();
      end
      endcase
    end
  end
  

endmodule

